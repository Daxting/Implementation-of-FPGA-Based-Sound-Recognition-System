`timescale 1ns / 10ps


module SignalPreAnalysis(
    input clk,
    input reset,
    input sound_input_Rready,
    input [15:0] sound_input,
    input log10_result_Wready,
    output reg sound_input_Wready,
    output reg [15:0] log10_result,
    output reg log10_result_Rready,
	output reg fftoff
    );
reg [2:0]NS, CS;
reg [15:0]hw_result[1023:0];
reg [15:0]fft_result[511:0];

parameter Initial = 3'd0, HWcal = 3'd1,SIwait = 3'd2, FFTcal = 3'd3, Melcal = 3'd4, Logtable = 3'd5, mfscout = 3'd6, waitram = 3'd7;

reg [9:0]hammingwindowAddr;
wire [15:0]HW_sel;
reg hammingwindowEnable;
reg SIread;
hamming_bank U0(.addra(hammingwindowAddr), .clka(clk), .douta(HW_sel), .ena(hammingwindowEnable));

reg[15:0] fft_input;
reg fft_s_axis_data_tvalid;
reg fft_s_axis_data_tlast;
wire fft_s_axis_data_tready;
wire fft_m_axis_data_tvalid;
wire fft_data_tvalid;
wire [15:0]fftout;
reg [9:0]fftinCount;
reg [8:0]fftoutCount;
reg fftfinish;

reg div_clk;
fft_modulus U1(clk, div_clk, reset, fft_input, fft_s_axis_data_tvalid, fft_s_axis_data_tlast,
fft_s_axis_data_tready, fft_m_axis_data_tvalid, fft_data_tvalid, fftout);

reg melbankEnable;
reg melfinish;
reg melcaldone;
reg [15:0] melout;
wire [15:0] mel_sel;
reg [14:0] melbankAddr;
reg [8:0]melcalCount;
reg [5:0]mfscoutCount;
melbank U2(.addra(melbankAddr), .clka(clk), .douta(mel_sel), .ena(melbankEnable));

reg logtablefinish;
reg [15:0] log10_cal;

// 50MHz clk
always@(posedge clk or negedge reset) begin
    if(!reset) begin
        div_clk <= 1'b0;
    end
    else begin
        div_clk <= !div_clk;
    end
end

//25MHz clk
reg divdiv_clk;
always@(posedge div_clk or negedge reset) begin
    if(!reset) begin
        divdiv_clk <= 1'b0;
    end
    else begin
        divdiv_clk <= !divdiv_clk;
    end
end

always@(posedge clk, negedge reset) begin
    if(!reset) begin
        CS <= 3'd0;
    end
    else begin
        CS <= NS;
    end
end

always@(*) begin
    case(CS)
        Initial: begin
            if(sound_input_Rready == 1'b1)
                NS = HWcal;
            else
                NS = Initial;
        end
        HWcal: begin
            if(sound_input_Rready == 1'b1 && SIread == 1'b1)
                NS = SIwait;
            else
                NS = HWcal;
        end
        SIwait: begin
            if(hammingwindowAddr == 10'd0)
                NS = FFTcal;
            else if(sound_input_Rready == 1'b1 && SIread == 1'b0)
                NS = HWcal;
            else
                NS = SIwait;
        end
        FFTcal: begin
            if(fftfinish == 1'b1)
                NS = Melcal;
            else
                NS = FFTcal;
        end
        Melcal: begin
            if(melcaldone == 1'b1)
                NS = Logtable;
            else
                NS = Melcal;
        end
        Logtable: begin
            if(logtablefinish == 1'b1)
                NS = mfscout;
            else
                NS = Logtable;
        end
        mfscout: begin
            if(log10_result_Wready == 1'b0)
                NS = waitram;
            else
                NS = mfscout;    
        end
        waitram: begin
            if(mfscoutCount == 6'd0 && log10_result_Wready == 1'b1)
                NS = Initial;
            else if(log10_result_Wready == 1'b1)
                NS = Melcal;
            else
                NS = waitram;
        end
        default: NS = Initial;
    endcase
end

always@(posedge clk or negedge reset) begin
    if(!reset) begin
        sound_input_Wready <= 1'b0;
        hammingwindowEnable <= 1'b0;
        fft_s_axis_data_tvalid <= 1'b0;
        fftoff <= 1'b0;
        melbankEnable <= 1'b0;
        melfinish <= 1'b0;
        log10_result_Rready <= 1'b0;
    end
    else begin
        case(CS)
            Initial: begin
                sound_input_Wready <= 1'b1;
                hammingwindowEnable <= 1'b1;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b0;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;
            end
            HWcal: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b1;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b0;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;   
            end
            SIwait: begin
                sound_input_Wready <= 1'b1;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b0;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;
            end
            FFTcal: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b1;
                fftoff <= 1'b0;
                melbankEnable <= 1'b1;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;
            end
            Melcal: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b1;
                melbankEnable <= 1'b1;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;
            end
            Logtable: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b1;
                melbankEnable <= 1'b0;
                melfinish <= 1'b1;
                log10_result_Rready <= 1'b0;
            end
            mfscout: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b1;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b1;
            end
            waitram: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b1;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b1;
            end
            default: begin
                sound_input_Wready <= 1'b0;
                hammingwindowEnable <= 1'b0;
                fft_s_axis_data_tvalid <= 1'b0;
                fftoff <= 1'b0;
                melbankEnable <= 1'b0;
                melfinish <= 1'b0;
                log10_result_Rready <= 1'b0;
            end
        endcase
    end
end

// hamming calculation
integer idx;
wire [31:0] partHWresult;
assign partHWresult = (sound_input[15] == 1'b1) ? {16'd65535, sound_input}*{16'd0, HW_sel}:
                                             {16'd0, sound_input}*{ 16'd0, HW_sel};
always@(posedge div_clk or negedge reset) begin
    if(!reset) begin
        hammingwindowAddr <= 10'd0;
        SIread <= 1'b0;
        for(idx=0; idx<1024; idx = idx + 1)begin
            hw_result[idx] <= 16'd0;
        end
    end
    else begin
        case(CS)
            HWcal: begin
                if(sound_input_Rready == 1'b1 && SIread <= 1'b0) begin
                    SIread <= 1'b1;
                    hammingwindowAddr <= hammingwindowAddr + 10'd1;
                    hw_result[hammingwindowAddr] <= {partHWresult[31], partHWresult[24:10]};
                end
                else begin
                    SIread <= 1'b0;
                    hammingwindowAddr <= hammingwindowAddr;
                    for(idx=0; idx<1024; idx = idx + 1)begin
                        hw_result[idx] <= hw_result[idx];
                    end
                end
            end
            SIwait: begin
               SIread <= 1'b0;
               hammingwindowAddr <= hammingwindowAddr;
               for(idx=0; idx<1024; idx = idx + 1)begin
                   hw_result[idx] <= hw_result[idx];
               end 
            end
            FFTcal: begin
                SIread <= 1'b0;
               hammingwindowAddr <= hammingwindowAddr;
               for(idx=0; idx<1024; idx = idx + 1)begin
                   hw_result[idx] <= hw_result[idx];
                end
            end
            default: begin
                SIread <= 1'b0;
                hammingwindowAddr <= 10'd0;
                for(idx=0; idx<1024; idx = idx + 1)begin
                    hw_result[idx] <= 16'd0;
                end
            end
        endcase
    end
end

// fftinput
always@(posedge div_clk or negedge reset) begin
    if(!reset) begin
        fft_input <= 16'd0;
        fftinCount <= 10'd0;
        fft_s_axis_data_tlast <= 1'b0;
    end
    else begin
        if(fft_s_axis_data_tready && fft_s_axis_data_tvalid) begin
            fft_input <= hw_result[fftinCount];
            fftinCount <= fftinCount + 10'd1;
            if(fftinCount == 10'd1023)
                fft_s_axis_data_tlast <= 1'b1;
            else
                fft_s_axis_data_tlast <= 1'b0;
        end
        else begin
            fft_input <= 16'd0;
            fftinCount <= 10'd0;
            fft_s_axis_data_tlast <= 1'b0;
        end
    end
end

//fft restoration
always@(posedge div_clk or negedge reset) begin
    if(!reset) begin
        for(idx=0; idx<512; idx = idx + 1)begin
            fft_result[idx] <= 16'd0;
        end
        fftoutCount <= 9'd0;
        fftfinish <= 1'b0;
    end
    else begin
        if(fft_m_axis_data_tvalid && fft_data_tvalid && fftoff == 1'b0) begin
            fft_result[fftoutCount] <= fftout;
            fftoutCount <= fftoutCount + 9'd1;
            if(fftoutCount == 9'd511)
                fftfinish <= 1'b1;
            else
                fftfinish <= 1'b0;
        end
        else begin
            for(idx=0; idx<512; idx = idx + 1)begin
                fft_result[idx] <= fft_result[idx];
            end
            fftoutCount <= 9'd0;
            fftfinish <= 1'b0; 
        end
    end
end

//melfilter
wire [31:0] partMelresult;
assign partMelresult = (fft_result[melcalCount][15] == 1'b1) ? {16'd65535, fft_result[melcalCount]}*{16'd0, mel_sel}:
                                                        {16'd0, fft_result[melcalCount]}*{ 16'd0, mel_sel};
always@(posedge divdiv_clk or negedge reset) begin
    if(!reset) begin
        melout <= 16'd0;
        melcalCount <= 9'd0;
        melbankAddr <= 15'd0;
        melcaldone <= 1'b0;
    end
    else begin
        case(CS)
            Melcal: begin
                if(fftoff == 1'b1) begin
                    melout <= melout + {partMelresult[31], partMelresult[24:10]};
                    melcalCount <= melcalCount + 9'd1;
                    melbankAddr <= melbankAddr + 15'd1;
                    if(melcalCount == 9'd511)
                        melcaldone <= 1'b1;
                    else
                        melcaldone <= 1'b0;
                end
                else begin
                    melout <= melout;
                    melcalCount <= melcalCount;
                    melbankAddr <= melbankAddr;
                    melcaldone <= 1'b0;
                end
            end
            Logtable: begin
                melout <= melout;
                melcalCount <= 9'd0;
                melbankAddr <= melbankAddr;
                melcaldone <= 1'b0;
            end
            mfscout: begin
                melout <= 16'd0;
                melcalCount <= 9'd0;
                melbankAddr <= melbankAddr;
                melcaldone <= 1'b0;
            end
            waitram: begin
                melout <= 16'd0;
                melcalCount <= 9'd0;
                melbankAddr <= melbankAddr;
                melcaldone <= 1'b0;
            end
            default: begin
                melout <= 16'd0;
                melcalCount <= 9'd0;
                melbankAddr <= 15'd0;
                melcaldone <= 1'b0;
            end
        endcase
    end
end

//logtable
always@(*)begin
    if(melfinish == 1'b1) begin
        case(melout[14:0])
            15'd1: log10_cal = 16'b1111001111110110;
            15'd2: log10_cal = 16'b1111010100101010;
            15'd3: log10_cal = 16'b1111010111011111;
            15'd4: log10_cal = 16'b1111011001011110;
            15'd5: log10_cal = 16'b1111011011000010;
            15'd6: log10_cal = 16'b1111011100010011;
            15'd7: log10_cal = 16'b1111011101010111;
            15'd8: log10_cal = 16'b1111011110010011;
            15'd9: log10_cal = 16'b1111011111000111;
            15'd10: log10_cal = 16'b1111011111110110;
            15'd11: log10_cal = 16'b1111100000100000;
            15'd12: log10_cal = 16'b1111100001000111;
            15'd13: log10_cal = 16'b1111100001101011;
            15'd14: log10_cal = 16'b1111100010001100;
            15'd15: log10_cal = 16'b1111100010101010;
            15'd16: log10_cal = 16'b1111100011000111;
            15'd17: log10_cal = 16'b1111100011100010;
            15'd18: log10_cal = 16'b1111100011111011;
            15'd19: log10_cal = 16'b1111100100010011;
            15'd20: log10_cal = 16'b1111100100101010;
            15'd21: log10_cal = 16'b1111100101000000;
            15'd22: log10_cal = 16'b1111100101010101;
            15'd23: log10_cal = 16'b1111100101101000;
            15'd24: log10_cal = 16'b1111100101111011;
            15'd25: log10_cal = 16'b1111100110001101;
            15'd26: log10_cal = 16'b1111100110011111;
            15'd27: log10_cal = 16'b1111100110110000;
            15'd28: log10_cal = 16'b1111100111000000;
            15'd29: log10_cal = 16'b1111100111001111;
            15'd30: log10_cal = 16'b1111100111011111;
            15'd31: log10_cal = 16'b1111100111101101;
            15'd32: log10_cal = 16'b1111100111111011;
            15'd33: log10_cal = 16'b1111101000001001;
            15'd34: log10_cal = 16'b1111101000010110;
            15'd35: log10_cal = 16'b1111101000100011;
            15'd36: log10_cal = 16'b1111101000110000;
            15'd37: log10_cal = 16'b1111101000111100;
            15'd38: log10_cal = 16'b1111101001001000;
            15'd39: log10_cal = 16'b1111101001010011;
            15'd40: log10_cal = 16'b1111101001011110;
            15'd41: log10_cal = 16'b1111101001101001;
            15'd42: log10_cal = 16'b1111101001110100;
            15'd43: log10_cal = 16'b1111101001111111;
            15'd44: log10_cal = 16'b1111101010001001;
            15'd45: log10_cal = 16'b1111101010010011;
            15'd46: log10_cal = 16'b1111101010011101;
            15'd47: log10_cal = 16'b1111101010100110;
            15'd48: log10_cal = 16'b1111101010110000;
            15'd49: log10_cal = 16'b1111101010111001;
            15'd50: log10_cal = 16'b1111101011000010;
            15'd51: log10_cal = 16'b1111101011001011;
            15'd52: log10_cal = 16'b1111101011010011;
            15'd53: log10_cal = 16'b1111101011011100;
            15'd54: log10_cal = 16'b1111101011100100;
            15'd55: log10_cal = 16'b1111101011101100;
            15'd56: log10_cal = 16'b1111101011110100;
            15'd57: log10_cal = 16'b1111101011111100;
            15'd58: log10_cal = 16'b1111101100000100;
            15'd59: log10_cal = 16'b1111101100001011;
            15'd60: log10_cal = 16'b1111101100010011;
            15'd61: log10_cal = 16'b1111101100011010;
            15'd62: log10_cal = 16'b1111101100100001;
            15'd63: log10_cal = 16'b1111101100101000;
            15'd64: log10_cal = 16'b1111101100101111;
            15'd65: log10_cal = 16'b1111101100110110;
            15'd66: log10_cal = 16'b1111101100111101;
            15'd67: log10_cal = 16'b1111101101000100;
            15'd68: log10_cal = 16'b1111101101001010;
            15'd69: log10_cal = 16'b1111101101010001;
            15'd70: log10_cal = 16'b1111101101010111;
            15'd71: log10_cal = 16'b1111101101011110;
            15'd72: log10_cal = 16'b1111101101100100;
            15'd73: log10_cal = 16'b1111101101101010;
            15'd74: log10_cal = 16'b1111101101110000;
            15'd75: log10_cal = 16'b1111101101110110;
            15'd76: log10_cal = 16'b1111101101111100;
            15'd77: log10_cal = 16'b1111101110000010;
            15'd78: log10_cal = 16'b1111101110000111;
            15'd79: log10_cal = 16'b1111101110001101;
            15'd80: log10_cal = 16'b1111101110010011;
            15'd81: log10_cal = 16'b1111101110011000;
            15'd82: log10_cal = 16'b1111101110011110;
            15'd83: log10_cal = 16'b1111101110100011;
            15'd84: log10_cal = 16'b1111101110101000;
            15'd85: log10_cal = 16'b1111101110101110;
            15'd86: log10_cal = 16'b1111101110110011;
            15'd87: log10_cal = 16'b1111101110111000;
            15'd88: log10_cal = 16'b1111101110111101;
            15'd89: log10_cal = 16'b1111101111000010;
            15'd90: log10_cal = 16'b1111101111000111;
            15'd91: log10_cal = 16'b1111101111001100;
            15'd92: log10_cal = 16'b1111101111010001;
            15'd93: log10_cal = 16'b1111101111010110;
            15'd94: log10_cal = 16'b1111101111011010;
            15'd95: log10_cal = 16'b1111101111011111;
            15'd96: log10_cal = 16'b1111101111100100;
            15'd97: log10_cal = 16'b1111101111101000;
            15'd98: log10_cal = 16'b1111101111101101;
            15'd99: log10_cal = 16'b1111101111110001;
            15'd100: log10_cal = 16'b1111101111110110;
            15'd101: log10_cal = 16'b1111101111111010;
            15'd102: log10_cal = 16'b1111101111111111;
            15'd103: log10_cal = 16'b1111110000000011;
            15'd104: log10_cal = 16'b1111110000000111;
            15'd105: log10_cal = 16'b1111110000001100;
            15'd106: log10_cal = 16'b1111110000010000;
            15'd107: log10_cal = 16'b1111110000010100;
            15'd108: log10_cal = 16'b1111110000011000;
            15'd109: log10_cal = 16'b1111110000011100;
            15'd110: log10_cal = 16'b1111110000100000;
            15'd111: log10_cal = 16'b1111110000100100;
            15'd112: log10_cal = 16'b1111110000101000;
            15'd113: log10_cal = 16'b1111110000101100;
            15'd114: log10_cal = 16'b1111110000110000;
            15'd115: log10_cal = 16'b1111110000110100;
            15'd116: log10_cal = 16'b1111110000111000;
            15'd117: log10_cal = 16'b1111110000111100;
            15'd118: log10_cal = 16'b1111110001000000;
            15'd119: log10_cal = 16'b1111110001000011;
            15'd120: log10_cal = 16'b1111110001000111;
            15'd121: log10_cal = 16'b1111110001001011;
            15'd122: log10_cal = 16'b1111110001001110;
            15'd123: log10_cal = 16'b1111110001010010;
            15'd124: log10_cal = 16'b1111110001010110;
            15'd125: log10_cal = 16'b1111110001011001;
            15'd126: log10_cal = 16'b1111110001011101;
            15'd127: log10_cal = 16'b1111110001100000;
            15'd128: log10_cal = 16'b1111110001100100;
            15'd129: log10_cal = 16'b1111110001100111;
            15'd130: log10_cal = 16'b1111110001101011;
            15'd131: log10_cal = 16'b1111110001101110;
            15'd132: log10_cal = 16'b1111110001110001;
            15'd133: log10_cal = 16'b1111110001110101;
            15'd134: log10_cal = 16'b1111110001111000;
            15'd135: log10_cal = 16'b1111110001111011;
            15'd136: log10_cal = 16'b1111110001111111;
            15'd137: log10_cal = 16'b1111110010000010;
            15'd138: log10_cal = 16'b1111110010000101;
            15'd139: log10_cal = 16'b1111110010001000;
            15'd140: log10_cal = 16'b1111110010001100;
            15'd141: log10_cal = 16'b1111110010001111;
            15'd142: log10_cal = 16'b1111110010010010;
            15'd143: log10_cal = 16'b1111110010010101;
            15'd144: log10_cal = 16'b1111110010011000;
            15'd145: log10_cal = 16'b1111110010011011;
            15'd146: log10_cal = 16'b1111110010011110;
            15'd147: log10_cal = 16'b1111110010100001;
            15'd148: log10_cal = 16'b1111110010100100;
            15'd149: log10_cal = 16'b1111110010100111;
            15'd150: log10_cal = 16'b1111110010101010;
            15'd151: log10_cal = 16'b1111110010101101;
            15'd152: log10_cal = 16'b1111110010110000;
            15'd153: log10_cal = 16'b1111110010110011;
            15'd154: log10_cal = 16'b1111110010110110;
            15'd155: log10_cal = 16'b1111110010111001;
            15'd156: log10_cal = 16'b1111110010111100;
            15'd157: log10_cal = 16'b1111110010111111;
            15'd158: log10_cal = 16'b1111110011000001;
            15'd159: log10_cal = 16'b1111110011000100;
            15'd160: log10_cal = 16'b1111110011000111;
            15'd161: log10_cal = 16'b1111110011001010;
            15'd162: log10_cal = 16'b1111110011001100;
            15'd163: log10_cal = 16'b1111110011001111;
            15'd164: log10_cal = 16'b1111110011010010;
            15'd165: log10_cal = 16'b1111110011010101;
            15'd166: log10_cal = 16'b1111110011010111;
            15'd167: log10_cal = 16'b1111110011011010;
            15'd168: log10_cal = 16'b1111110011011101;
            15'd169: log10_cal = 16'b1111110011011111;
            15'd170: log10_cal = 16'b1111110011100010;
            15'd171: log10_cal = 16'b1111110011100101;
            15'd172: log10_cal = 16'b1111110011100111;
            15'd173: log10_cal = 16'b1111110011101010;
            15'd174: log10_cal = 16'b1111110011101100;
            15'd175: log10_cal = 16'b1111110011101111;
            15'd176: log10_cal = 16'b1111110011110001;
            15'd177: log10_cal = 16'b1111110011110100;
            15'd178: log10_cal = 16'b1111110011110110;
            15'd179: log10_cal = 16'b1111110011111001;
            15'd180: log10_cal = 16'b1111110011111011;
            15'd181: log10_cal = 16'b1111110011111110;
            15'd182: log10_cal = 16'b1111110100000000;
            15'd183: log10_cal = 16'b1111110100000011;
            15'd184: log10_cal = 16'b1111110100000101;
            15'd185: log10_cal = 16'b1111110100001000;
            15'd186: log10_cal = 16'b1111110100001010;
            15'd187: log10_cal = 16'b1111110100001100;
            15'd188: log10_cal = 16'b1111110100001111;
            15'd189: log10_cal = 16'b1111110100010001;
            15'd190: log10_cal = 16'b1111110100010011;
            15'd191: log10_cal = 16'b1111110100010110;
            15'd192: log10_cal = 16'b1111110100011000;
            15'd193: log10_cal = 16'b1111110100011010;
            15'd194: log10_cal = 16'b1111110100011101;
            15'd195: log10_cal = 16'b1111110100011111;
            15'd196: log10_cal = 16'b1111110100100001;
            15'd197: log10_cal = 16'b1111110100100011;
            15'd198: log10_cal = 16'b1111110100100110;
            15'd199: log10_cal = 16'b1111110100101000;
            15'd200: log10_cal = 16'b1111110100101010;
            15'd201: log10_cal = 16'b1111110100101100;
            15'd202: log10_cal = 16'b1111110100101111;
            15'd203: log10_cal = 16'b1111110100110001;
            15'd204: log10_cal = 16'b1111110100110011;
            15'd205: log10_cal = 16'b1111110100110101;
            15'd206: log10_cal = 16'b1111110100110111;
            15'd207: log10_cal = 16'b1111110100111010;
            15'd208: log10_cal = 16'b1111110100111100;
            15'd209: log10_cal = 16'b1111110100111110;
            15'd210: log10_cal = 16'b1111110101000000;
            15'd211: log10_cal = 16'b1111110101000010;
            15'd212: log10_cal = 16'b1111110101000100;
            15'd213: log10_cal = 16'b1111110101000110;
            15'd214: log10_cal = 16'b1111110101001000;
            15'd215: log10_cal = 16'b1111110101001010;
            15'd216: log10_cal = 16'b1111110101001100;
            15'd217: log10_cal = 16'b1111110101001110;
            15'd218: log10_cal = 16'b1111110101010001;
            15'd219: log10_cal = 16'b1111110101010011;
            15'd220: log10_cal = 16'b1111110101010101;
            15'd221: log10_cal = 16'b1111110101010111;
            15'd222: log10_cal = 16'b1111110101011001;
            15'd223: log10_cal = 16'b1111110101011011;
            15'd224: log10_cal = 16'b1111110101011101;
            15'd225: log10_cal = 16'b1111110101011111;
            15'd226: log10_cal = 16'b1111110101100001;
            15'd227: log10_cal = 16'b1111110101100011;
            15'd228: log10_cal = 16'b1111110101100100;
            15'd229: log10_cal = 16'b1111110101100110;
            15'd230: log10_cal = 16'b1111110101101000;
            15'd231: log10_cal = 16'b1111110101101010;
            15'd232: log10_cal = 16'b1111110101101100;
            15'd233: log10_cal = 16'b1111110101101110;
            15'd234: log10_cal = 16'b1111110101110000;
            15'd235: log10_cal = 16'b1111110101110010;
            15'd236: log10_cal = 16'b1111110101110100;
            15'd237: log10_cal = 16'b1111110101110110;
            15'd238: log10_cal = 16'b1111110101111000;
            15'd239: log10_cal = 16'b1111110101111001;
            15'd240: log10_cal = 16'b1111110101111011;
            15'd241: log10_cal = 16'b1111110101111101;
            15'd242: log10_cal = 16'b1111110101111111;
            15'd243: log10_cal = 16'b1111110110000001;
            15'd244: log10_cal = 16'b1111110110000011;
            15'd245: log10_cal = 16'b1111110110000100;
            15'd246: log10_cal = 16'b1111110110000110;
            15'd247: log10_cal = 16'b1111110110001000;
            15'd248: log10_cal = 16'b1111110110001010;
            15'd249: log10_cal = 16'b1111110110001100;
            15'd250: log10_cal = 16'b1111110110001101;
            15'd251: log10_cal = 16'b1111110110001111;
            15'd252: log10_cal = 16'b1111110110010001;
            15'd253: log10_cal = 16'b1111110110010011;
            15'd254: log10_cal = 16'b1111110110010101;
            15'd255: log10_cal = 16'b1111110110010110;
            15'd256: log10_cal = 16'b1111110110011000;
            15'd257: log10_cal = 16'b1111110110011010;
            15'd258: log10_cal = 16'b1111110110011011;
            15'd259: log10_cal = 16'b1111110110011101;
            15'd260: log10_cal = 16'b1111110110011111;
            15'd261: log10_cal = 16'b1111110110100001;
            15'd262: log10_cal = 16'b1111110110100010;
            15'd263: log10_cal = 16'b1111110110100100;
            15'd264: log10_cal = 16'b1111110110100110;
            15'd265: log10_cal = 16'b1111110110100111;
            15'd266: log10_cal = 16'b1111110110101001;
            15'd267: log10_cal = 16'b1111110110101011;
            15'd268: log10_cal = 16'b1111110110101100;
            15'd269: log10_cal = 16'b1111110110101110;
            15'd270: log10_cal = 16'b1111110110110000;
            15'd271: log10_cal = 16'b1111110110110001;
            15'd272: log10_cal = 16'b1111110110110011;
            15'd273: log10_cal = 16'b1111110110110101;
            15'd274: log10_cal = 16'b1111110110110110;
            15'd275: log10_cal = 16'b1111110110111000;
            15'd276: log10_cal = 16'b1111110110111001;
            15'd277: log10_cal = 16'b1111110110111011;
            15'd278: log10_cal = 16'b1111110110111101;
            15'd279: log10_cal = 16'b1111110110111110;
            15'd280: log10_cal = 16'b1111110111000000;
            15'd281: log10_cal = 16'b1111110111000001;
            15'd282: log10_cal = 16'b1111110111000011;
            15'd283: log10_cal = 16'b1111110111000101;
            15'd284: log10_cal = 16'b1111110111000110;
            15'd285: log10_cal = 16'b1111110111001000;
            15'd286: log10_cal = 16'b1111110111001001;
            15'd287: log10_cal = 16'b1111110111001011;
            15'd288: log10_cal = 16'b1111110111001100;
            15'd289: log10_cal = 16'b1111110111001110;
            15'd290: log10_cal = 16'b1111110111001111;
            15'd291: log10_cal = 16'b1111110111010001;
            15'd292: log10_cal = 16'b1111110111010011;
            15'd293: log10_cal = 16'b1111110111010100;
            15'd294: log10_cal = 16'b1111110111010110;
            15'd295: log10_cal = 16'b1111110111010111;
            15'd296: log10_cal = 16'b1111110111011001;
            15'd297: log10_cal = 16'b1111110111011010;
            15'd298: log10_cal = 16'b1111110111011100;
            15'd299: log10_cal = 16'b1111110111011101;
            15'd300: log10_cal = 16'b1111110111011111;
            15'd301: log10_cal = 16'b1111110111100000;
            15'd302: log10_cal = 16'b1111110111100001;
            15'd303: log10_cal = 16'b1111110111100011;
            15'd304: log10_cal = 16'b1111110111100100;
            15'd305: log10_cal = 16'b1111110111100110;
            15'd306: log10_cal = 16'b1111110111100111;
            15'd307: log10_cal = 16'b1111110111101001;
            15'd308: log10_cal = 16'b1111110111101010;
            15'd309: log10_cal = 16'b1111110111101100;
            15'd310: log10_cal = 16'b1111110111101101;
            15'd311: log10_cal = 16'b1111110111101111;
            15'd312: log10_cal = 16'b1111110111110000;
            15'd313: log10_cal = 16'b1111110111110001;
            15'd314: log10_cal = 16'b1111110111110011;
            15'd315: log10_cal = 16'b1111110111110100;
            15'd316: log10_cal = 16'b1111110111110110;
            15'd317: log10_cal = 16'b1111110111110111;
            15'd318: log10_cal = 16'b1111110111111000;
            15'd319: log10_cal = 16'b1111110111111010;
            15'd320: log10_cal = 16'b1111110111111011;
            15'd321: log10_cal = 16'b1111110111111101;
            15'd322: log10_cal = 16'b1111110111111110;
            15'd323: log10_cal = 16'b1111110111111111;
            15'd324: log10_cal = 16'b1111111000000001;
            15'd325: log10_cal = 16'b1111111000000010;
            15'd326: log10_cal = 16'b1111111000000011;
            15'd327: log10_cal = 16'b1111111000000101;
            15'd328: log10_cal = 16'b1111111000000110;
            15'd329: log10_cal = 16'b1111111000001000;
            15'd330: log10_cal = 16'b1111111000001001;
            15'd331: log10_cal = 16'b1111111000001010;
            15'd332: log10_cal = 16'b1111111000001100;
            15'd333: log10_cal = 16'b1111111000001101;
            15'd334: log10_cal = 16'b1111111000001110;
            15'd335: log10_cal = 16'b1111111000010000;
            15'd336: log10_cal = 16'b1111111000010001;
            15'd337: log10_cal = 16'b1111111000010010;
            15'd338: log10_cal = 16'b1111111000010100;
            15'd339: log10_cal = 16'b1111111000010101;
            15'd340: log10_cal = 16'b1111111000010110;
            15'd341: log10_cal = 16'b1111111000010111;
            15'd342: log10_cal = 16'b1111111000011001;
            15'd343: log10_cal = 16'b1111111000011010;
            15'd344: log10_cal = 16'b1111111000011011;
            15'd345: log10_cal = 16'b1111111000011101;
            15'd346: log10_cal = 16'b1111111000011110;
            15'd347: log10_cal = 16'b1111111000011111;
            15'd348: log10_cal = 16'b1111111000100001;
            15'd349: log10_cal = 16'b1111111000100010;
            15'd350: log10_cal = 16'b1111111000100011;
            15'd351: log10_cal = 16'b1111111000100100;
            15'd352: log10_cal = 16'b1111111000100110;
            15'd353: log10_cal = 16'b1111111000100111;
            15'd354: log10_cal = 16'b1111111000101000;
            15'd355: log10_cal = 16'b1111111000101001;
            15'd356: log10_cal = 16'b1111111000101011;
            15'd357: log10_cal = 16'b1111111000101100;
            15'd358: log10_cal = 16'b1111111000101101;
            15'd359: log10_cal = 16'b1111111000101110;
            15'd360: log10_cal = 16'b1111111000110000;
            15'd361: log10_cal = 16'b1111111000110001;
            15'd362: log10_cal = 16'b1111111000110010;
            15'd363: log10_cal = 16'b1111111000110011;
            15'd364: log10_cal = 16'b1111111000110101;
            15'd365: log10_cal = 16'b1111111000110110;
            15'd366: log10_cal = 16'b1111111000110111;
            15'd367: log10_cal = 16'b1111111000111000;
            15'd368: log10_cal = 16'b1111111000111001;
            15'd369: log10_cal = 16'b1111111000111011;
            15'd370: log10_cal = 16'b1111111000111100;
            15'd371: log10_cal = 16'b1111111000111101;
            15'd372: log10_cal = 16'b1111111000111110;
            15'd373: log10_cal = 16'b1111111000111111;
            15'd374: log10_cal = 16'b1111111001000001;
            15'd375: log10_cal = 16'b1111111001000010;
            15'd376: log10_cal = 16'b1111111001000011;
            15'd377: log10_cal = 16'b1111111001000100;
            15'd378: log10_cal = 16'b1111111001000101;
            15'd379: log10_cal = 16'b1111111001000110;
            15'd380: log10_cal = 16'b1111111001001000;
            15'd381: log10_cal = 16'b1111111001001001;
            15'd382: log10_cal = 16'b1111111001001010;
            15'd383: log10_cal = 16'b1111111001001011;
            15'd384: log10_cal = 16'b1111111001001100;
            15'd385: log10_cal = 16'b1111111001001101;
            15'd386: log10_cal = 16'b1111111001001111;
            15'd387: log10_cal = 16'b1111111001010000;
            15'd388: log10_cal = 16'b1111111001010001;
            15'd389: log10_cal = 16'b1111111001010010;
            15'd390: log10_cal = 16'b1111111001010011;
            15'd391: log10_cal = 16'b1111111001010100;
            15'd392: log10_cal = 16'b1111111001010101;
            15'd393: log10_cal = 16'b1111111001010111;
            15'd394: log10_cal = 16'b1111111001011000;
            15'd395: log10_cal = 16'b1111111001011001;
            15'd396: log10_cal = 16'b1111111001011010;
            15'd397: log10_cal = 16'b1111111001011011;
            15'd398: log10_cal = 16'b1111111001011100;
            15'd399: log10_cal = 16'b1111111001011101;
            15'd400: log10_cal = 16'b1111111001011110;
            15'd401: log10_cal = 16'b1111111001100000;
            15'd402: log10_cal = 16'b1111111001100001;
            15'd403: log10_cal = 16'b1111111001100010;
            15'd404: log10_cal = 16'b1111111001100011;
            15'd405: log10_cal = 16'b1111111001100100;
            15'd406: log10_cal = 16'b1111111001100101;
            15'd407: log10_cal = 16'b1111111001100110;
            15'd408: log10_cal = 16'b1111111001100111;
            15'd409: log10_cal = 16'b1111111001101000;
            15'd410: log10_cal = 16'b1111111001101001;
            15'd411: log10_cal = 16'b1111111001101011;
            15'd412: log10_cal = 16'b1111111001101100;
            15'd413: log10_cal = 16'b1111111001101101;
            15'd414: log10_cal = 16'b1111111001101110;
            15'd415: log10_cal = 16'b1111111001101111;
            15'd416: log10_cal = 16'b1111111001110000;
            15'd417: log10_cal = 16'b1111111001110001;
            15'd418: log10_cal = 16'b1111111001110010;
            15'd419: log10_cal = 16'b1111111001110011;
            15'd420: log10_cal = 16'b1111111001110100;
            15'd421: log10_cal = 16'b1111111001110101;
            15'd422: log10_cal = 16'b1111111001110110;
            15'd423: log10_cal = 16'b1111111001110111;
            15'd424: log10_cal = 16'b1111111001111000;
            15'd425: log10_cal = 16'b1111111001111001;
            15'd426: log10_cal = 16'b1111111001111010;
            15'd427: log10_cal = 16'b1111111001111100;
            15'd428: log10_cal = 16'b1111111001111101;
            15'd429: log10_cal = 16'b1111111001111110;
            15'd430: log10_cal = 16'b1111111001111111;
            15'd431: log10_cal = 16'b1111111010000000;
            15'd432: log10_cal = 16'b1111111010000001;
            15'd433: log10_cal = 16'b1111111010000010;
            15'd434: log10_cal = 16'b1111111010000011;
            15'd435: log10_cal = 16'b1111111010000100;
            15'd436: log10_cal = 16'b1111111010000101;
            15'd437: log10_cal = 16'b1111111010000110;
            15'd438: log10_cal = 16'b1111111010000111;
            15'd439: log10_cal = 16'b1111111010001000;
            15'd440: log10_cal = 16'b1111111010001001;
            15'd441: log10_cal = 16'b1111111010001010;
            15'd442: log10_cal = 16'b1111111010001011;
            15'd443: log10_cal = 16'b1111111010001100;
            15'd444: log10_cal = 16'b1111111010001101;
            15'd445: log10_cal = 16'b1111111010001110;
            15'd446: log10_cal = 16'b1111111010001111;
            15'd447: log10_cal = 16'b1111111010010000;
            15'd448: log10_cal = 16'b1111111010010001;
            15'd449: log10_cal = 16'b1111111010010010;
            15'd450: log10_cal = 16'b1111111010010011;
            15'd451: log10_cal = 16'b1111111010010100;
            15'd452: log10_cal = 16'b1111111010010101;
            15'd453: log10_cal = 16'b1111111010010110;
            15'd454: log10_cal = 16'b1111111010010111;
            15'd455: log10_cal = 16'b1111111010011000;
            15'd456: log10_cal = 16'b1111111010011001;
            15'd457: log10_cal = 16'b1111111010011010;
            15'd458: log10_cal = 16'b1111111010011011;
            15'd459: log10_cal = 16'b1111111010011100;
            15'd460: log10_cal = 16'b1111111010011101;
            15'd461: log10_cal = 16'b1111111010011110;
            15'd462: log10_cal = 16'b1111111010011111;
            15'd463: log10_cal = 16'b1111111010100000;
            15'd464: log10_cal = 16'b1111111010100000;
            15'd465: log10_cal = 16'b1111111010100001;
            15'd466: log10_cal = 16'b1111111010100010;
            15'd467: log10_cal = 16'b1111111010100011;
            15'd468: log10_cal = 16'b1111111010100100;
            15'd469: log10_cal = 16'b1111111010100101;
            15'd470: log10_cal = 16'b1111111010100110;
            15'd471: log10_cal = 16'b1111111010100111;
            15'd472: log10_cal = 16'b1111111010101000;
            15'd473: log10_cal = 16'b1111111010101001;
            15'd474: log10_cal = 16'b1111111010101010;
            15'd475: log10_cal = 16'b1111111010101011;
            15'd476: log10_cal = 16'b1111111010101100;
            15'd477: log10_cal = 16'b1111111010101101;
            15'd478: log10_cal = 16'b1111111010101110;
            15'd479: log10_cal = 16'b1111111010101111;
            15'd480: log10_cal = 16'b1111111010110000;
            15'd481: log10_cal = 16'b1111111010110000;
            15'd482: log10_cal = 16'b1111111010110001;
            15'd483: log10_cal = 16'b1111111010110010;
            15'd484: log10_cal = 16'b1111111010110011;
            15'd485: log10_cal = 16'b1111111010110100;
            15'd486: log10_cal = 16'b1111111010110101;
            15'd487: log10_cal = 16'b1111111010110110;
            15'd488: log10_cal = 16'b1111111010110111;
            15'd489: log10_cal = 16'b1111111010111000;
            15'd490: log10_cal = 16'b1111111010111001;
            15'd491: log10_cal = 16'b1111111010111010;
            15'd492: log10_cal = 16'b1111111010111011;
            15'd493: log10_cal = 16'b1111111010111011;
            15'd494: log10_cal = 16'b1111111010111100;
            15'd495: log10_cal = 16'b1111111010111101;
            15'd496: log10_cal = 16'b1111111010111110;
            15'd497: log10_cal = 16'b1111111010111111;
            15'd498: log10_cal = 16'b1111111011000000;
            15'd499: log10_cal = 16'b1111111011000001;
            15'd500: log10_cal = 16'b1111111011000010;
            15'd501: log10_cal = 16'b1111111011000011;
            15'd502: log10_cal = 16'b1111111011000011;
            15'd503: log10_cal = 16'b1111111011000100;
            15'd504: log10_cal = 16'b1111111011000101;
            15'd505: log10_cal = 16'b1111111011000110;
            15'd506: log10_cal = 16'b1111111011000111;
            15'd507: log10_cal = 16'b1111111011001000;
            15'd508: log10_cal = 16'b1111111011001001;
            15'd509: log10_cal = 16'b1111111011001010;
            15'd510: log10_cal = 16'b1111111011001011;
            15'd511: log10_cal = 16'b1111111011001011;
            15'd512: log10_cal = 16'b1111111011001100;
            15'd513: log10_cal = 16'b1111111011001101;
            15'd514: log10_cal = 16'b1111111011001110;
            15'd515: log10_cal = 16'b1111111011001111;
            15'd516: log10_cal = 16'b1111111011010000;
            15'd517: log10_cal = 16'b1111111011010001;
            15'd518: log10_cal = 16'b1111111011010001;
            15'd519: log10_cal = 16'b1111111011010010;
            15'd520: log10_cal = 16'b1111111011010011;
            15'd521: log10_cal = 16'b1111111011010100;
            15'd522: log10_cal = 16'b1111111011010101;
            15'd523: log10_cal = 16'b1111111011010110;
            15'd524: log10_cal = 16'b1111111011010111;
            15'd525: log10_cal = 16'b1111111011010111;
            15'd526: log10_cal = 16'b1111111011011000;
            15'd527: log10_cal = 16'b1111111011011001;
            15'd528: log10_cal = 16'b1111111011011010;
            15'd529: log10_cal = 16'b1111111011011011;
            15'd530: log10_cal = 16'b1111111011011100;
            15'd531: log10_cal = 16'b1111111011011100;
            15'd532: log10_cal = 16'b1111111011011101;
            15'd533: log10_cal = 16'b1111111011011110;
            15'd534: log10_cal = 16'b1111111011011111;
            15'd535: log10_cal = 16'b1111111011100000;
            15'd536: log10_cal = 16'b1111111011100001;
            15'd537: log10_cal = 16'b1111111011100001;
            15'd538: log10_cal = 16'b1111111011100010;
            15'd539: log10_cal = 16'b1111111011100011;
            15'd540: log10_cal = 16'b1111111011100100;
            15'd541: log10_cal = 16'b1111111011100101;
            15'd542: log10_cal = 16'b1111111011100110;
            15'd543: log10_cal = 16'b1111111011100110;
            15'd544: log10_cal = 16'b1111111011100111;
            15'd545: log10_cal = 16'b1111111011101000;
            15'd546: log10_cal = 16'b1111111011101001;
            15'd547: log10_cal = 16'b1111111011101010;
            15'd548: log10_cal = 16'b1111111011101010;
            15'd549: log10_cal = 16'b1111111011101011;
            15'd550: log10_cal = 16'b1111111011101100;
            15'd551: log10_cal = 16'b1111111011101101;
            15'd552: log10_cal = 16'b1111111011101110;
            15'd553: log10_cal = 16'b1111111011101111;
            15'd554: log10_cal = 16'b1111111011101111;
            15'd555: log10_cal = 16'b1111111011110000;
            15'd556: log10_cal = 16'b1111111011110001;
            15'd557: log10_cal = 16'b1111111011110010;
            15'd558: log10_cal = 16'b1111111011110011;
            15'd559: log10_cal = 16'b1111111011110011;
            15'd560: log10_cal = 16'b1111111011110100;
            15'd561: log10_cal = 16'b1111111011110101;
            15'd562: log10_cal = 16'b1111111011110110;
            15'd563: log10_cal = 16'b1111111011110110;
            15'd564: log10_cal = 16'b1111111011110111;
            15'd565: log10_cal = 16'b1111111011111000;
            15'd566: log10_cal = 16'b1111111011111001;
            15'd567: log10_cal = 16'b1111111011111010;
            15'd568: log10_cal = 16'b1111111011111010;
            15'd569: log10_cal = 16'b1111111011111011;
            15'd570: log10_cal = 16'b1111111011111100;
            15'd571: log10_cal = 16'b1111111011111101;
            15'd572: log10_cal = 16'b1111111011111110;
            15'd573: log10_cal = 16'b1111111011111110;
            15'd574: log10_cal = 16'b1111111011111111;
            15'd575: log10_cal = 16'b1111111100000000;
            15'd576: log10_cal = 16'b1111111100000001;
            15'd577: log10_cal = 16'b1111111100000001;
            15'd578: log10_cal = 16'b1111111100000010;
            15'd579: log10_cal = 16'b1111111100000011;
            15'd580: log10_cal = 16'b1111111100000100;
            15'd581: log10_cal = 16'b1111111100000100;
            15'd582: log10_cal = 16'b1111111100000101;
            15'd583: log10_cal = 16'b1111111100000110;
            15'd584: log10_cal = 16'b1111111100000111;
            15'd585: log10_cal = 16'b1111111100001000;
            15'd586: log10_cal = 16'b1111111100001000;
            15'd587: log10_cal = 16'b1111111100001001;
            15'd588: log10_cal = 16'b1111111100001010;
            15'd589: log10_cal = 16'b1111111100001011;
            15'd590: log10_cal = 16'b1111111100001011;
            15'd591: log10_cal = 16'b1111111100001100;
            15'd592: log10_cal = 16'b1111111100001101;
            15'd593: log10_cal = 16'b1111111100001110;
            15'd594: log10_cal = 16'b1111111100001110;
            15'd595: log10_cal = 16'b1111111100001111;
            15'd596: log10_cal = 16'b1111111100010000;
            15'd597: log10_cal = 16'b1111111100010001;
            15'd598: log10_cal = 16'b1111111100010001;
            15'd599: log10_cal = 16'b1111111100010010;
            15'd600: log10_cal = 16'b1111111100010011;
            15'd601: log10_cal = 16'b1111111100010100;
            15'd602: log10_cal = 16'b1111111100010100;
            15'd603: log10_cal = 16'b1111111100010101;
            15'd604: log10_cal = 16'b1111111100010110;
            15'd605: log10_cal = 16'b1111111100010110;
            15'd606: log10_cal = 16'b1111111100010111;
            15'd607: log10_cal = 16'b1111111100011000;
            15'd608: log10_cal = 16'b1111111100011001;
            15'd609: log10_cal = 16'b1111111100011001;
            15'd610: log10_cal = 16'b1111111100011010;
            15'd611: log10_cal = 16'b1111111100011011;
            15'd612: log10_cal = 16'b1111111100011100;
            15'd613: log10_cal = 16'b1111111100011100;
            15'd614: log10_cal = 16'b1111111100011101;
            15'd615: log10_cal = 16'b1111111100011110;
            15'd616: log10_cal = 16'b1111111100011110;
            15'd617: log10_cal = 16'b1111111100011111;
            15'd618: log10_cal = 16'b1111111100100000;
            15'd619: log10_cal = 16'b1111111100100001;
            15'd620: log10_cal = 16'b1111111100100001;
            15'd621: log10_cal = 16'b1111111100100010;
            15'd622: log10_cal = 16'b1111111100100011;
            15'd623: log10_cal = 16'b1111111100100100;
            15'd624: log10_cal = 16'b1111111100100100;
            15'd625: log10_cal = 16'b1111111100100101;
            15'd626: log10_cal = 16'b1111111100100110;
            15'd627: log10_cal = 16'b1111111100100110;
            15'd628: log10_cal = 16'b1111111100100111;
            15'd629: log10_cal = 16'b1111111100101000;
            15'd630: log10_cal = 16'b1111111100101000;
            15'd631: log10_cal = 16'b1111111100101001;
            15'd632: log10_cal = 16'b1111111100101010;
            15'd633: log10_cal = 16'b1111111100101011;
            15'd634: log10_cal = 16'b1111111100101011;
            15'd635: log10_cal = 16'b1111111100101100;
            15'd636: log10_cal = 16'b1111111100101101;
            15'd637: log10_cal = 16'b1111111100101101;
            15'd638: log10_cal = 16'b1111111100101110;
            15'd639: log10_cal = 16'b1111111100101111;
            15'd640: log10_cal = 16'b1111111100101111;
            15'd641: log10_cal = 16'b1111111100110000;
            15'd642: log10_cal = 16'b1111111100110001;
            15'd643: log10_cal = 16'b1111111100110010;
            15'd644: log10_cal = 16'b1111111100110010;
            15'd645: log10_cal = 16'b1111111100110011;
            15'd646: log10_cal = 16'b1111111100110100;
            15'd647: log10_cal = 16'b1111111100110100;
            15'd648: log10_cal = 16'b1111111100110101;
            15'd649: log10_cal = 16'b1111111100110110;
            15'd650: log10_cal = 16'b1111111100110110;
            15'd651: log10_cal = 16'b1111111100110111;
            15'd652: log10_cal = 16'b1111111100111000;
            15'd653: log10_cal = 16'b1111111100111000;
            15'd654: log10_cal = 16'b1111111100111001;
            15'd655: log10_cal = 16'b1111111100111010;
            15'd656: log10_cal = 16'b1111111100111010;
            15'd657: log10_cal = 16'b1111111100111011;
            15'd658: log10_cal = 16'b1111111100111100;
            15'd659: log10_cal = 16'b1111111100111100;
            15'd660: log10_cal = 16'b1111111100111101;
            15'd661: log10_cal = 16'b1111111100111110;
            15'd662: log10_cal = 16'b1111111100111111;
            15'd663: log10_cal = 16'b1111111100111111;
            15'd664: log10_cal = 16'b1111111101000000;
            15'd665: log10_cal = 16'b1111111101000001;
            15'd666: log10_cal = 16'b1111111101000001;
            15'd667: log10_cal = 16'b1111111101000010;
            15'd668: log10_cal = 16'b1111111101000011;
            15'd669: log10_cal = 16'b1111111101000011;
            15'd670: log10_cal = 16'b1111111101000100;
            15'd671: log10_cal = 16'b1111111101000101;
            15'd672: log10_cal = 16'b1111111101000101;
            15'd673: log10_cal = 16'b1111111101000110;
            15'd674: log10_cal = 16'b1111111101000111;
            15'd675: log10_cal = 16'b1111111101000111;
            15'd676: log10_cal = 16'b1111111101001000;
            15'd677: log10_cal = 16'b1111111101001000;
            15'd678: log10_cal = 16'b1111111101001001;
            15'd679: log10_cal = 16'b1111111101001010;
            15'd680: log10_cal = 16'b1111111101001010;
            15'd681: log10_cal = 16'b1111111101001011;
            15'd682: log10_cal = 16'b1111111101001100;
            15'd683: log10_cal = 16'b1111111101001100;
            15'd684: log10_cal = 16'b1111111101001101;
            15'd685: log10_cal = 16'b1111111101001110;
            15'd686: log10_cal = 16'b1111111101001110;
            15'd687: log10_cal = 16'b1111111101001111;
            15'd688: log10_cal = 16'b1111111101010000;
            15'd689: log10_cal = 16'b1111111101010000;
            15'd690: log10_cal = 16'b1111111101010001;
            15'd691: log10_cal = 16'b1111111101010010;
            15'd692: log10_cal = 16'b1111111101010010;
            15'd693: log10_cal = 16'b1111111101010011;
            15'd694: log10_cal = 16'b1111111101010100;
            15'd695: log10_cal = 16'b1111111101010100;
            15'd696: log10_cal = 16'b1111111101010101;
            15'd697: log10_cal = 16'b1111111101010101;
            15'd698: log10_cal = 16'b1111111101010110;
            15'd699: log10_cal = 16'b1111111101010111;
            15'd700: log10_cal = 16'b1111111101010111;
            15'd701: log10_cal = 16'b1111111101011000;
            15'd702: log10_cal = 16'b1111111101011001;
            15'd703: log10_cal = 16'b1111111101011001;
            15'd704: log10_cal = 16'b1111111101011010;
            15'd705: log10_cal = 16'b1111111101011010;
            15'd706: log10_cal = 16'b1111111101011011;
            15'd707: log10_cal = 16'b1111111101011100;
            15'd708: log10_cal = 16'b1111111101011100;
            15'd709: log10_cal = 16'b1111111101011101;
            15'd710: log10_cal = 16'b1111111101011110;
            15'd711: log10_cal = 16'b1111111101011110;
            15'd712: log10_cal = 16'b1111111101011111;
            15'd713: log10_cal = 16'b1111111101100000;
            15'd714: log10_cal = 16'b1111111101100000;
            15'd715: log10_cal = 16'b1111111101100001;
            15'd716: log10_cal = 16'b1111111101100001;
            15'd717: log10_cal = 16'b1111111101100010;
            15'd718: log10_cal = 16'b1111111101100011;
            15'd719: log10_cal = 16'b1111111101100011;
            15'd720: log10_cal = 16'b1111111101100100;
            15'd721: log10_cal = 16'b1111111101100100;
            15'd722: log10_cal = 16'b1111111101100101;
            15'd723: log10_cal = 16'b1111111101100110;
            15'd724: log10_cal = 16'b1111111101100110;
            15'd725: log10_cal = 16'b1111111101100111;
            15'd726: log10_cal = 16'b1111111101101000;
            15'd727: log10_cal = 16'b1111111101101000;
            15'd728: log10_cal = 16'b1111111101101001;
            15'd729: log10_cal = 16'b1111111101101001;
            15'd730: log10_cal = 16'b1111111101101010;
            15'd731: log10_cal = 16'b1111111101101011;
            15'd732: log10_cal = 16'b1111111101101011;
            15'd733: log10_cal = 16'b1111111101101100;
            15'd734: log10_cal = 16'b1111111101101100;
            15'd735: log10_cal = 16'b1111111101101101;
            15'd736: log10_cal = 16'b1111111101101110;
            15'd737: log10_cal = 16'b1111111101101110;
            15'd738: log10_cal = 16'b1111111101101111;
            15'd739: log10_cal = 16'b1111111101101111;
            15'd740: log10_cal = 16'b1111111101110000;
            15'd741: log10_cal = 16'b1111111101110001;
            15'd742: log10_cal = 16'b1111111101110001;
            15'd743: log10_cal = 16'b1111111101110010;
            15'd744: log10_cal = 16'b1111111101110010;
            15'd745: log10_cal = 16'b1111111101110011;
            15'd746: log10_cal = 16'b1111111101110100;
            15'd747: log10_cal = 16'b1111111101110100;
            15'd748: log10_cal = 16'b1111111101110101;
            15'd749: log10_cal = 16'b1111111101110101;
            15'd750: log10_cal = 16'b1111111101110110;
            15'd751: log10_cal = 16'b1111111101110111;
            15'd752: log10_cal = 16'b1111111101110111;
            15'd753: log10_cal = 16'b1111111101111000;
            15'd754: log10_cal = 16'b1111111101111000;
            15'd755: log10_cal = 16'b1111111101111001;
            15'd756: log10_cal = 16'b1111111101111010;
            15'd757: log10_cal = 16'b1111111101111010;
            15'd758: log10_cal = 16'b1111111101111011;
            15'd759: log10_cal = 16'b1111111101111011;
            15'd760: log10_cal = 16'b1111111101111100;
            15'd761: log10_cal = 16'b1111111101111100;
            15'd762: log10_cal = 16'b1111111101111101;
            15'd763: log10_cal = 16'b1111111101111110;
            15'd764: log10_cal = 16'b1111111101111110;
            15'd765: log10_cal = 16'b1111111101111111;
            15'd766: log10_cal = 16'b1111111101111111;
            15'd767: log10_cal = 16'b1111111110000000;
            15'd768: log10_cal = 16'b1111111110000001;
            15'd769: log10_cal = 16'b1111111110000001;
            15'd770: log10_cal = 16'b1111111110000010;
            15'd771: log10_cal = 16'b1111111110000010;
            15'd772: log10_cal = 16'b1111111110000011;
            15'd773: log10_cal = 16'b1111111110000011;
            15'd774: log10_cal = 16'b1111111110000100;
            15'd775: log10_cal = 16'b1111111110000101;
            15'd776: log10_cal = 16'b1111111110000101;
            15'd777: log10_cal = 16'b1111111110000110;
            15'd778: log10_cal = 16'b1111111110000110;
            15'd779: log10_cal = 16'b1111111110000111;
            15'd780: log10_cal = 16'b1111111110000111;
            15'd781: log10_cal = 16'b1111111110001000;
            15'd782: log10_cal = 16'b1111111110001001;
            15'd783: log10_cal = 16'b1111111110001001;
            15'd784: log10_cal = 16'b1111111110001010;
            15'd785: log10_cal = 16'b1111111110001010;
            15'd786: log10_cal = 16'b1111111110001011;
            15'd787: log10_cal = 16'b1111111110001011;
            15'd788: log10_cal = 16'b1111111110001100;
            15'd789: log10_cal = 16'b1111111110001101;
            15'd790: log10_cal = 16'b1111111110001101;
            15'd791: log10_cal = 16'b1111111110001110;
            15'd792: log10_cal = 16'b1111111110001110;
            15'd793: log10_cal = 16'b1111111110001111;
            15'd794: log10_cal = 16'b1111111110001111;
            15'd795: log10_cal = 16'b1111111110010000;
            15'd796: log10_cal = 16'b1111111110010000;
            15'd797: log10_cal = 16'b1111111110010001;
            15'd798: log10_cal = 16'b1111111110010010;
            15'd799: log10_cal = 16'b1111111110010010;
            15'd800: log10_cal = 16'b1111111110010011;
            15'd801: log10_cal = 16'b1111111110010011;
            15'd802: log10_cal = 16'b1111111110010100;
            15'd803: log10_cal = 16'b1111111110010100;
            15'd804: log10_cal = 16'b1111111110010101;
            15'd805: log10_cal = 16'b1111111110010101;
            15'd806: log10_cal = 16'b1111111110010110;
            15'd807: log10_cal = 16'b1111111110010111;
            15'd808: log10_cal = 16'b1111111110010111;
            15'd809: log10_cal = 16'b1111111110011000;
            15'd810: log10_cal = 16'b1111111110011000;
            15'd811: log10_cal = 16'b1111111110011001;
            15'd812: log10_cal = 16'b1111111110011001;
            15'd813: log10_cal = 16'b1111111110011010;
            15'd814: log10_cal = 16'b1111111110011010;
            15'd815: log10_cal = 16'b1111111110011011;
            15'd816: log10_cal = 16'b1111111110011100;
            15'd817: log10_cal = 16'b1111111110011100;
            15'd818: log10_cal = 16'b1111111110011101;
            15'd819: log10_cal = 16'b1111111110011101;
            15'd820: log10_cal = 16'b1111111110011110;
            15'd821: log10_cal = 16'b1111111110011110;
            15'd822: log10_cal = 16'b1111111110011111;
            15'd823: log10_cal = 16'b1111111110011111;
            15'd824: log10_cal = 16'b1111111110100000;
            15'd825: log10_cal = 16'b1111111110100000;
            15'd826: log10_cal = 16'b1111111110100001;
            15'd827: log10_cal = 16'b1111111110100001;
            15'd828: log10_cal = 16'b1111111110100010;
            15'd829: log10_cal = 16'b1111111110100011;
            15'd830: log10_cal = 16'b1111111110100011;
            15'd831: log10_cal = 16'b1111111110100100;
            15'd832: log10_cal = 16'b1111111110100100;
            15'd833: log10_cal = 16'b1111111110100101;
            15'd834: log10_cal = 16'b1111111110100101;
            15'd835: log10_cal = 16'b1111111110100110;
            15'd836: log10_cal = 16'b1111111110100110;
            15'd837: log10_cal = 16'b1111111110100111;
            15'd838: log10_cal = 16'b1111111110100111;
            15'd839: log10_cal = 16'b1111111110101000;
            15'd840: log10_cal = 16'b1111111110101000;
            15'd841: log10_cal = 16'b1111111110101001;
            15'd842: log10_cal = 16'b1111111110101001;
            15'd843: log10_cal = 16'b1111111110101010;
            15'd844: log10_cal = 16'b1111111110101011;
            15'd845: log10_cal = 16'b1111111110101011;
            15'd846: log10_cal = 16'b1111111110101100;
            15'd847: log10_cal = 16'b1111111110101100;
            15'd848: log10_cal = 16'b1111111110101101;
            15'd849: log10_cal = 16'b1111111110101101;
            15'd850: log10_cal = 16'b1111111110101110;
            15'd851: log10_cal = 16'b1111111110101110;
            15'd852: log10_cal = 16'b1111111110101111;
            15'd853: log10_cal = 16'b1111111110101111;
            15'd854: log10_cal = 16'b1111111110110000;
            15'd855: log10_cal = 16'b1111111110110000;
            15'd856: log10_cal = 16'b1111111110110001;
            15'd857: log10_cal = 16'b1111111110110001;
            15'd858: log10_cal = 16'b1111111110110010;
            15'd859: log10_cal = 16'b1111111110110010;
            15'd860: log10_cal = 16'b1111111110110011;
            15'd861: log10_cal = 16'b1111111110110011;
            15'd862: log10_cal = 16'b1111111110110100;
            15'd863: log10_cal = 16'b1111111110110100;
            15'd864: log10_cal = 16'b1111111110110101;
            15'd865: log10_cal = 16'b1111111110110101;
            15'd866: log10_cal = 16'b1111111110110110;
            15'd867: log10_cal = 16'b1111111110110110;
            15'd868: log10_cal = 16'b1111111110110111;
            15'd869: log10_cal = 16'b1111111110111000;
            15'd870: log10_cal = 16'b1111111110111000;
            15'd871: log10_cal = 16'b1111111110111001;
            15'd872: log10_cal = 16'b1111111110111001;
            15'd873: log10_cal = 16'b1111111110111010;
            15'd874: log10_cal = 16'b1111111110111010;
            15'd875: log10_cal = 16'b1111111110111011;
            15'd876: log10_cal = 16'b1111111110111011;
            15'd877: log10_cal = 16'b1111111110111100;
            15'd878: log10_cal = 16'b1111111110111100;
            15'd879: log10_cal = 16'b1111111110111101;
            15'd880: log10_cal = 16'b1111111110111101;
            15'd881: log10_cal = 16'b1111111110111110;
            15'd882: log10_cal = 16'b1111111110111110;
            15'd883: log10_cal = 16'b1111111110111111;
            15'd884: log10_cal = 16'b1111111110111111;
            15'd885: log10_cal = 16'b1111111111000000;
            15'd886: log10_cal = 16'b1111111111000000;
            15'd887: log10_cal = 16'b1111111111000001;
            15'd888: log10_cal = 16'b1111111111000001;
            15'd889: log10_cal = 16'b1111111111000010;
            15'd890: log10_cal = 16'b1111111111000010;
            15'd891: log10_cal = 16'b1111111111000011;
            15'd892: log10_cal = 16'b1111111111000011;
            15'd893: log10_cal = 16'b1111111111000100;
            15'd894: log10_cal = 16'b1111111111000100;
            15'd895: log10_cal = 16'b1111111111000101;
            15'd896: log10_cal = 16'b1111111111000101;
            15'd897: log10_cal = 16'b1111111111000110;
            15'd898: log10_cal = 16'b1111111111000110;
            15'd899: log10_cal = 16'b1111111111000111;
            15'd900: log10_cal = 16'b1111111111000111;
            15'd901: log10_cal = 16'b1111111111001000;
            15'd902: log10_cal = 16'b1111111111001000;
            15'd903: log10_cal = 16'b1111111111001001;
            15'd904: log10_cal = 16'b1111111111001001;
            15'd905: log10_cal = 16'b1111111111001010;
            15'd906: log10_cal = 16'b1111111111001010;
            15'd907: log10_cal = 16'b1111111111001011;
            15'd908: log10_cal = 16'b1111111111001011;
            15'd909: log10_cal = 16'b1111111111001100;
            15'd910: log10_cal = 16'b1111111111001100;
            15'd911: log10_cal = 16'b1111111111001100;
            15'd912: log10_cal = 16'b1111111111001101;
            15'd913: log10_cal = 16'b1111111111001101;
            15'd914: log10_cal = 16'b1111111111001110;
            15'd915: log10_cal = 16'b1111111111001110;
            15'd916: log10_cal = 16'b1111111111001111;
            15'd917: log10_cal = 16'b1111111111001111;
            15'd918: log10_cal = 16'b1111111111010000;
            15'd919: log10_cal = 16'b1111111111010000;
            15'd920: log10_cal = 16'b1111111111010001;
            15'd921: log10_cal = 16'b1111111111010001;
            15'd922: log10_cal = 16'b1111111111010010;
            15'd923: log10_cal = 16'b1111111111010010;
            15'd924: log10_cal = 16'b1111111111010011;
            15'd925: log10_cal = 16'b1111111111010011;
            15'd926: log10_cal = 16'b1111111111010100;
            15'd927: log10_cal = 16'b1111111111010100;
            15'd928: log10_cal = 16'b1111111111010101;
            15'd929: log10_cal = 16'b1111111111010101;
            15'd930: log10_cal = 16'b1111111111010110;
            15'd931: log10_cal = 16'b1111111111010110;
            15'd932: log10_cal = 16'b1111111111010111;
            15'd933: log10_cal = 16'b1111111111010111;
            15'd934: log10_cal = 16'b1111111111011000;
            15'd935: log10_cal = 16'b1111111111011000;
            15'd936: log10_cal = 16'b1111111111011001;
            15'd937: log10_cal = 16'b1111111111011001;
            15'd938: log10_cal = 16'b1111111111011001;
            15'd939: log10_cal = 16'b1111111111011010;
            15'd940: log10_cal = 16'b1111111111011010;
            15'd941: log10_cal = 16'b1111111111011011;
            15'd942: log10_cal = 16'b1111111111011011;
            15'd943: log10_cal = 16'b1111111111011100;
            15'd944: log10_cal = 16'b1111111111011100;
            15'd945: log10_cal = 16'b1111111111011101;
            15'd946: log10_cal = 16'b1111111111011101;
            15'd947: log10_cal = 16'b1111111111011110;
            15'd948: log10_cal = 16'b1111111111011110;
            15'd949: log10_cal = 16'b1111111111011111;
            15'd950: log10_cal = 16'b1111111111011111;
            15'd951: log10_cal = 16'b1111111111100000;
            15'd952: log10_cal = 16'b1111111111100000;
            15'd953: log10_cal = 16'b1111111111100001;
            15'd954: log10_cal = 16'b1111111111100001;
            15'd955: log10_cal = 16'b1111111111100001;
            15'd956: log10_cal = 16'b1111111111100010;
            15'd957: log10_cal = 16'b1111111111100010;
            15'd958: log10_cal = 16'b1111111111100011;
            15'd959: log10_cal = 16'b1111111111100011;
            15'd960: log10_cal = 16'b1111111111100100;
            15'd961: log10_cal = 16'b1111111111100100;
            15'd962: log10_cal = 16'b1111111111100101;
            15'd963: log10_cal = 16'b1111111111100101;
            15'd964: log10_cal = 16'b1111111111100110;
            15'd965: log10_cal = 16'b1111111111100110;
            15'd966: log10_cal = 16'b1111111111100111;
            15'd967: log10_cal = 16'b1111111111100111;
            15'd968: log10_cal = 16'b1111111111100111;
            15'd969: log10_cal = 16'b1111111111101000;
            15'd970: log10_cal = 16'b1111111111101000;
            15'd971: log10_cal = 16'b1111111111101001;
            15'd972: log10_cal = 16'b1111111111101001;
            15'd973: log10_cal = 16'b1111111111101010;
            15'd974: log10_cal = 16'b1111111111101010;
            15'd975: log10_cal = 16'b1111111111101011;
            15'd976: log10_cal = 16'b1111111111101011;
            15'd977: log10_cal = 16'b1111111111101100;
            15'd978: log10_cal = 16'b1111111111101100;
            15'd979: log10_cal = 16'b1111111111101101;
            15'd980: log10_cal = 16'b1111111111101101;
            15'd981: log10_cal = 16'b1111111111101101;
            15'd982: log10_cal = 16'b1111111111101110;
            15'd983: log10_cal = 16'b1111111111101110;
            15'd984: log10_cal = 16'b1111111111101111;
            15'd985: log10_cal = 16'b1111111111101111;
            15'd986: log10_cal = 16'b1111111111110000;
            15'd987: log10_cal = 16'b1111111111110000;
            15'd988: log10_cal = 16'b1111111111110001;
            15'd989: log10_cal = 16'b1111111111110001;
            15'd990: log10_cal = 16'b1111111111110001;
            15'd991: log10_cal = 16'b1111111111110010;
            15'd992: log10_cal = 16'b1111111111110010;
            15'd993: log10_cal = 16'b1111111111110011;
            15'd994: log10_cal = 16'b1111111111110011;
            15'd995: log10_cal = 16'b1111111111110100;
            15'd996: log10_cal = 16'b1111111111110100;
            15'd997: log10_cal = 16'b1111111111110101;
            15'd998: log10_cal = 16'b1111111111110101;
            15'd999: log10_cal = 16'b1111111111110110;
            15'd1000: log10_cal = 16'b1111111111110110;
            15'd1001: log10_cal = 16'b1111111111110110;
            15'd1002: log10_cal = 16'b1111111111110111;
            15'd1003: log10_cal = 16'b1111111111110111;
            15'd1004: log10_cal = 16'b1111111111111000;
            15'd1005: log10_cal = 16'b1111111111111000;
            15'd1006: log10_cal = 16'b1111111111111001;
            15'd1007: log10_cal = 16'b1111111111111001;
            15'd1008: log10_cal = 16'b1111111111111001;
            15'd1009: log10_cal = 16'b1111111111111010;
            15'd1010: log10_cal = 16'b1111111111111010;
            15'd1011: log10_cal = 16'b1111111111111011;
            15'd1012: log10_cal = 16'b1111111111111011;
            15'd1013: log10_cal = 16'b1111111111111100;
            15'd1014: log10_cal = 16'b1111111111111100;
            15'd1015: log10_cal = 16'b1111111111111101;
            15'd1016: log10_cal = 16'b1111111111111101;
            15'd1017: log10_cal = 16'b1111111111111101;
            15'd1018: log10_cal = 16'b1111111111111110;
            15'd1019: log10_cal = 16'b1111111111111110;
            15'd1020: log10_cal = 16'b1111111111111111;
            15'd1021: log10_cal = 16'b1111111111111111;
            15'd1022: log10_cal = 16'b1000000000000000;
            15'd1023: log10_cal = 16'b1000000000000000;
            15'd1024: log10_cal = 16'b0000000000000000;
            15'd1025: log10_cal = 16'b0000000000000000;
            15'd1026: log10_cal = 16'b0000000000000000;
            15'd1027: log10_cal = 16'b0000000000000001;
            15'd1028: log10_cal = 16'b0000000000000001;
            15'd1029: log10_cal = 16'b0000000000000010;
            15'd1030: log10_cal = 16'b0000000000000010;
            15'd1031: log10_cal = 16'b0000000000000011;
            15'd1032: log10_cal = 16'b0000000000000011;
            15'd1033: log10_cal = 16'b0000000000000011;
            15'd1034: log10_cal = 16'b0000000000000100;
            15'd1035: log10_cal = 16'b0000000000000100;
            15'd1036: log10_cal = 16'b0000000000000101;
            15'd1037: log10_cal = 16'b0000000000000101;
            15'd1038: log10_cal = 16'b0000000000000110;
            15'd1039: log10_cal = 16'b0000000000000110;
            15'd1040: log10_cal = 16'b0000000000000110;
            15'd1041: log10_cal = 16'b0000000000000111;
            15'd1042: log10_cal = 16'b0000000000000111;
            15'd1043: log10_cal = 16'b0000000000001000;
            15'd1044: log10_cal = 16'b0000000000001000;
            15'd1045: log10_cal = 16'b0000000000001001;
            15'd1046: log10_cal = 16'b0000000000001001;
            15'd1047: log10_cal = 16'b0000000000001001;
            15'd1048: log10_cal = 16'b0000000000001010;
            15'd1049: log10_cal = 16'b0000000000001010;
            15'd1050: log10_cal = 16'b0000000000001011;
            15'd1051: log10_cal = 16'b0000000000001011;
            15'd1052: log10_cal = 16'b0000000000001011;
            15'd1053: log10_cal = 16'b0000000000001100;
            15'd1054: log10_cal = 16'b0000000000001100;
            15'd1055: log10_cal = 16'b0000000000001101;
            15'd1056: log10_cal = 16'b0000000000001101;
            15'd1057: log10_cal = 16'b0000000000001110;
            15'd1058: log10_cal = 16'b0000000000001110;
            15'd1059: log10_cal = 16'b0000000000001110;
            15'd1060: log10_cal = 16'b0000000000001111;
            15'd1061: log10_cal = 16'b0000000000001111;
            15'd1062: log10_cal = 16'b0000000000010000;
            15'd1063: log10_cal = 16'b0000000000010000;
            15'd1064: log10_cal = 16'b0000000000010001;
            15'd1065: log10_cal = 16'b0000000000010001;
            15'd1066: log10_cal = 16'b0000000000010001;
            15'd1067: log10_cal = 16'b0000000000010010;
            15'd1068: log10_cal = 16'b0000000000010010;
            15'd1069: log10_cal = 16'b0000000000010011;
            15'd1070: log10_cal = 16'b0000000000010011;
            15'd1071: log10_cal = 16'b0000000000010011;
            15'd1072: log10_cal = 16'b0000000000010100;
            15'd1073: log10_cal = 16'b0000000000010100;
            15'd1074: log10_cal = 16'b0000000000010101;
            15'd1075: log10_cal = 16'b0000000000010101;
            15'd1076: log10_cal = 16'b0000000000010110;
            15'd1077: log10_cal = 16'b0000000000010110;
            15'd1078: log10_cal = 16'b0000000000010110;
            15'd1079: log10_cal = 16'b0000000000010111;
            15'd1080: log10_cal = 16'b0000000000010111;
            15'd1081: log10_cal = 16'b0000000000011000;
            15'd1082: log10_cal = 16'b0000000000011000;
            15'd1083: log10_cal = 16'b0000000000011000;
            15'd1084: log10_cal = 16'b0000000000011001;
            15'd1085: log10_cal = 16'b0000000000011001;
            15'd1086: log10_cal = 16'b0000000000011010;
            15'd1087: log10_cal = 16'b0000000000011010;
            15'd1088: log10_cal = 16'b0000000000011010;
            15'd1089: log10_cal = 16'b0000000000011011;
            15'd1090: log10_cal = 16'b0000000000011011;
            15'd1091: log10_cal = 16'b0000000000011100;
            15'd1092: log10_cal = 16'b0000000000011100;
            15'd1093: log10_cal = 16'b0000000000011100;
            15'd1094: log10_cal = 16'b0000000000011101;
            15'd1095: log10_cal = 16'b0000000000011101;
            15'd1096: log10_cal = 16'b0000000000011110;
            15'd1097: log10_cal = 16'b0000000000011110;
            15'd1098: log10_cal = 16'b0000000000011111;
            15'd1099: log10_cal = 16'b0000000000011111;
            15'd1100: log10_cal = 16'b0000000000011111;
            15'd1101: log10_cal = 16'b0000000000100000;
            15'd1102: log10_cal = 16'b0000000000100000;
            15'd1103: log10_cal = 16'b0000000000100001;
            15'd1104: log10_cal = 16'b0000000000100001;
            15'd1105: log10_cal = 16'b0000000000100001;
            15'd1106: log10_cal = 16'b0000000000100010;
            15'd1107: log10_cal = 16'b0000000000100010;
            15'd1108: log10_cal = 16'b0000000000100011;
            15'd1109: log10_cal = 16'b0000000000100011;
            15'd1110: log10_cal = 16'b0000000000100011;
            15'd1111: log10_cal = 16'b0000000000100100;
            15'd1112: log10_cal = 16'b0000000000100100;
            15'd1113: log10_cal = 16'b0000000000100101;
            15'd1114: log10_cal = 16'b0000000000100101;
            15'd1115: log10_cal = 16'b0000000000100101;
            15'd1116: log10_cal = 16'b0000000000100110;
            15'd1117: log10_cal = 16'b0000000000100110;
            15'd1118: log10_cal = 16'b0000000000100111;
            15'd1119: log10_cal = 16'b0000000000100111;
            15'd1120: log10_cal = 16'b0000000000100111;
            15'd1121: log10_cal = 16'b0000000000101000;
            15'd1122: log10_cal = 16'b0000000000101000;
            15'd1123: log10_cal = 16'b0000000000101001;
            15'd1124: log10_cal = 16'b0000000000101001;
            15'd1125: log10_cal = 16'b0000000000101001;
            15'd1126: log10_cal = 16'b0000000000101010;
            15'd1127: log10_cal = 16'b0000000000101010;
            15'd1128: log10_cal = 16'b0000000000101011;
            15'd1129: log10_cal = 16'b0000000000101011;
            15'd1130: log10_cal = 16'b0000000000101011;
            15'd1131: log10_cal = 16'b0000000000101100;
            15'd1132: log10_cal = 16'b0000000000101100;
            15'd1133: log10_cal = 16'b0000000000101100;
            15'd1134: log10_cal = 16'b0000000000101101;
            15'd1135: log10_cal = 16'b0000000000101101;
            15'd1136: log10_cal = 16'b0000000000101110;
            15'd1137: log10_cal = 16'b0000000000101110;
            15'd1138: log10_cal = 16'b0000000000101110;
            15'd1139: log10_cal = 16'b0000000000101111;
            15'd1140: log10_cal = 16'b0000000000101111;
            15'd1141: log10_cal = 16'b0000000000110000;
            15'd1142: log10_cal = 16'b0000000000110000;
            15'd1143: log10_cal = 16'b0000000000110000;
            15'd1144: log10_cal = 16'b0000000000110001;
            15'd1145: log10_cal = 16'b0000000000110001;
            15'd1146: log10_cal = 16'b0000000000110010;
            15'd1147: log10_cal = 16'b0000000000110010;
            15'd1148: log10_cal = 16'b0000000000110010;
            15'd1149: log10_cal = 16'b0000000000110011;
            15'd1150: log10_cal = 16'b0000000000110011;
            15'd1151: log10_cal = 16'b0000000000110011;
            15'd1152: log10_cal = 16'b0000000000110100;
            15'd1153: log10_cal = 16'b0000000000110100;
            15'd1154: log10_cal = 16'b0000000000110101;
            15'd1155: log10_cal = 16'b0000000000110101;
            15'd1156: log10_cal = 16'b0000000000110101;
            15'd1157: log10_cal = 16'b0000000000110110;
            15'd1158: log10_cal = 16'b0000000000110110;
            15'd1159: log10_cal = 16'b0000000000110111;
            15'd1160: log10_cal = 16'b0000000000110111;
            15'd1161: log10_cal = 16'b0000000000110111;
            15'd1162: log10_cal = 16'b0000000000111000;
            15'd1163: log10_cal = 16'b0000000000111000;
            15'd1164: log10_cal = 16'b0000000000111000;
            15'd1165: log10_cal = 16'b0000000000111001;
            15'd1166: log10_cal = 16'b0000000000111001;
            15'd1167: log10_cal = 16'b0000000000111010;
            15'd1168: log10_cal = 16'b0000000000111010;
            15'd1169: log10_cal = 16'b0000000000111010;
            15'd1170: log10_cal = 16'b0000000000111011;
            15'd1171: log10_cal = 16'b0000000000111011;
            15'd1172: log10_cal = 16'b0000000000111100;
            15'd1173: log10_cal = 16'b0000000000111100;
            15'd1174: log10_cal = 16'b0000000000111100;
            15'd1175: log10_cal = 16'b0000000000111101;
            15'd1176: log10_cal = 16'b0000000000111101;
            15'd1177: log10_cal = 16'b0000000000111101;
            15'd1178: log10_cal = 16'b0000000000111110;
            15'd1179: log10_cal = 16'b0000000000111110;
            15'd1180: log10_cal = 16'b0000000000111111;
            15'd1181: log10_cal = 16'b0000000000111111;
            15'd1182: log10_cal = 16'b0000000000111111;
            15'd1183: log10_cal = 16'b0000000001000000;
            15'd1184: log10_cal = 16'b0000000001000000;
            15'd1185: log10_cal = 16'b0000000001000000;
            15'd1186: log10_cal = 16'b0000000001000001;
            15'd1187: log10_cal = 16'b0000000001000001;
            15'd1188: log10_cal = 16'b0000000001000010;
            15'd1189: log10_cal = 16'b0000000001000010;
            15'd1190: log10_cal = 16'b0000000001000010;
            15'd1191: log10_cal = 16'b0000000001000011;
            15'd1192: log10_cal = 16'b0000000001000011;
            15'd1193: log10_cal = 16'b0000000001000011;
            15'd1194: log10_cal = 16'b0000000001000100;
            15'd1195: log10_cal = 16'b0000000001000100;
            15'd1196: log10_cal = 16'b0000000001000101;
            15'd1197: log10_cal = 16'b0000000001000101;
            15'd1198: log10_cal = 16'b0000000001000101;
            15'd1199: log10_cal = 16'b0000000001000110;
            15'd1200: log10_cal = 16'b0000000001000110;
            15'd1201: log10_cal = 16'b0000000001000110;
            15'd1202: log10_cal = 16'b0000000001000111;
            15'd1203: log10_cal = 16'b0000000001000111;
            15'd1204: log10_cal = 16'b0000000001001000;
            15'd1205: log10_cal = 16'b0000000001001000;
            15'd1206: log10_cal = 16'b0000000001001000;
            15'd1207: log10_cal = 16'b0000000001001001;
            15'd1208: log10_cal = 16'b0000000001001001;
            15'd1209: log10_cal = 16'b0000000001001001;
            15'd1210: log10_cal = 16'b0000000001001010;
            15'd1211: log10_cal = 16'b0000000001001010;
            15'd1212: log10_cal = 16'b0000000001001010;
            15'd1213: log10_cal = 16'b0000000001001011;
            15'd1214: log10_cal = 16'b0000000001001011;
            15'd1215: log10_cal = 16'b0000000001001100;
            15'd1216: log10_cal = 16'b0000000001001100;
            15'd1217: log10_cal = 16'b0000000001001100;
            15'd1218: log10_cal = 16'b0000000001001101;
            15'd1219: log10_cal = 16'b0000000001001101;
            15'd1220: log10_cal = 16'b0000000001001101;
            15'd1221: log10_cal = 16'b0000000001001110;
            15'd1222: log10_cal = 16'b0000000001001110;
            15'd1223: log10_cal = 16'b0000000001001110;
            15'd1224: log10_cal = 16'b0000000001001111;
            15'd1225: log10_cal = 16'b0000000001001111;
            15'd1226: log10_cal = 16'b0000000001010000;
            15'd1227: log10_cal = 16'b0000000001010000;
            15'd1228: log10_cal = 16'b0000000001010000;
            15'd1229: log10_cal = 16'b0000000001010001;
            15'd1230: log10_cal = 16'b0000000001010001;
            15'd1231: log10_cal = 16'b0000000001010001;
            15'd1232: log10_cal = 16'b0000000001010010;
            15'd1233: log10_cal = 16'b0000000001010010;
            15'd1234: log10_cal = 16'b0000000001010010;
            15'd1235: log10_cal = 16'b0000000001010011;
            15'd1236: log10_cal = 16'b0000000001010011;
            15'd1237: log10_cal = 16'b0000000001010100;
            15'd1238: log10_cal = 16'b0000000001010100;
            15'd1239: log10_cal = 16'b0000000001010100;
            15'd1240: log10_cal = 16'b0000000001010101;
            15'd1241: log10_cal = 16'b0000000001010101;
            15'd1242: log10_cal = 16'b0000000001010101;
            15'd1243: log10_cal = 16'b0000000001010110;
            15'd1244: log10_cal = 16'b0000000001010110;
            15'd1245: log10_cal = 16'b0000000001010110;
            15'd1246: log10_cal = 16'b0000000001010111;
            15'd1247: log10_cal = 16'b0000000001010111;
            15'd1248: log10_cal = 16'b0000000001010111;
            15'd1249: log10_cal = 16'b0000000001011000;
            15'd1250: log10_cal = 16'b0000000001011000;
            15'd1251: log10_cal = 16'b0000000001011001;
            15'd1252: log10_cal = 16'b0000000001011001;
            15'd1253: log10_cal = 16'b0000000001011001;
            15'd1254: log10_cal = 16'b0000000001011010;
            15'd1255: log10_cal = 16'b0000000001011010;
            15'd1256: log10_cal = 16'b0000000001011010;
            15'd1257: log10_cal = 16'b0000000001011011;
            15'd1258: log10_cal = 16'b0000000001011011;
            15'd1259: log10_cal = 16'b0000000001011011;
            15'd1260: log10_cal = 16'b0000000001011100;
            15'd1261: log10_cal = 16'b0000000001011100;
            15'd1262: log10_cal = 16'b0000000001011100;
            15'd1263: log10_cal = 16'b0000000001011101;
            15'd1264: log10_cal = 16'b0000000001011101;
            15'd1265: log10_cal = 16'b0000000001011101;
            15'd1266: log10_cal = 16'b0000000001011110;
            15'd1267: log10_cal = 16'b0000000001011110;
            15'd1268: log10_cal = 16'b0000000001011111;
            15'd1269: log10_cal = 16'b0000000001011111;
            15'd1270: log10_cal = 16'b0000000001011111;
            15'd1271: log10_cal = 16'b0000000001100000;
            15'd1272: log10_cal = 16'b0000000001100000;
            15'd1273: log10_cal = 16'b0000000001100000;
            15'd1274: log10_cal = 16'b0000000001100001;
            15'd1275: log10_cal = 16'b0000000001100001;
            15'd1276: log10_cal = 16'b0000000001100001;
            15'd1277: log10_cal = 16'b0000000001100010;
            15'd1278: log10_cal = 16'b0000000001100010;
            15'd1279: log10_cal = 16'b0000000001100010;
            15'd1280: log10_cal = 16'b0000000001100011;
            15'd1281: log10_cal = 16'b0000000001100011;
            15'd1282: log10_cal = 16'b0000000001100011;
            15'd1283: log10_cal = 16'b0000000001100100;
            15'd1284: log10_cal = 16'b0000000001100100;
            15'd1285: log10_cal = 16'b0000000001100100;
            15'd1286: log10_cal = 16'b0000000001100101;
            15'd1287: log10_cal = 16'b0000000001100101;
            15'd1288: log10_cal = 16'b0000000001100110;
            15'd1289: log10_cal = 16'b0000000001100110;
            15'd1290: log10_cal = 16'b0000000001100110;
            15'd1291: log10_cal = 16'b0000000001100111;
            15'd1292: log10_cal = 16'b0000000001100111;
            15'd1293: log10_cal = 16'b0000000001100111;
            15'd1294: log10_cal = 16'b0000000001101000;
            15'd1295: log10_cal = 16'b0000000001101000;
            15'd1296: log10_cal = 16'b0000000001101000;
            15'd1297: log10_cal = 16'b0000000001101001;
            15'd1298: log10_cal = 16'b0000000001101001;
            15'd1299: log10_cal = 16'b0000000001101001;
            15'd1300: log10_cal = 16'b0000000001101010;
            15'd1301: log10_cal = 16'b0000000001101010;
            15'd1302: log10_cal = 16'b0000000001101010;
            15'd1303: log10_cal = 16'b0000000001101011;
            15'd1304: log10_cal = 16'b0000000001101011;
            15'd1305: log10_cal = 16'b0000000001101011;
            15'd1306: log10_cal = 16'b0000000001101100;
            15'd1307: log10_cal = 16'b0000000001101100;
            15'd1308: log10_cal = 16'b0000000001101100;
            15'd1309: log10_cal = 16'b0000000001101101;
            15'd1310: log10_cal = 16'b0000000001101101;
            15'd1311: log10_cal = 16'b0000000001101101;
            15'd1312: log10_cal = 16'b0000000001101110;
            15'd1313: log10_cal = 16'b0000000001101110;
            15'd1314: log10_cal = 16'b0000000001101110;
            15'd1315: log10_cal = 16'b0000000001101111;
            15'd1316: log10_cal = 16'b0000000001101111;
            15'd1317: log10_cal = 16'b0000000001101111;
            15'd1318: log10_cal = 16'b0000000001110000;
            15'd1319: log10_cal = 16'b0000000001110000;
            15'd1320: log10_cal = 16'b0000000001110000;
            15'd1321: log10_cal = 16'b0000000001110001;
            15'd1322: log10_cal = 16'b0000000001110001;
            15'd1323: log10_cal = 16'b0000000001110001;
            15'd1324: log10_cal = 16'b0000000001110010;
            15'd1325: log10_cal = 16'b0000000001110010;
            15'd1326: log10_cal = 16'b0000000001110010;
            15'd1327: log10_cal = 16'b0000000001110011;
            15'd1328: log10_cal = 16'b0000000001110011;
            15'd1329: log10_cal = 16'b0000000001110011;
            15'd1330: log10_cal = 16'b0000000001110100;
            15'd1331: log10_cal = 16'b0000000001110100;
            15'd1332: log10_cal = 16'b0000000001110100;
            15'd1333: log10_cal = 16'b0000000001110101;
            15'd1334: log10_cal = 16'b0000000001110101;
            15'd1335: log10_cal = 16'b0000000001110101;
            15'd1336: log10_cal = 16'b0000000001110110;
            15'd1337: log10_cal = 16'b0000000001110110;
            15'd1338: log10_cal = 16'b0000000001110110;
            15'd1339: log10_cal = 16'b0000000001110111;
            15'd1340: log10_cal = 16'b0000000001110111;
            15'd1341: log10_cal = 16'b0000000001110111;
            15'd1342: log10_cal = 16'b0000000001111000;
            15'd1343: log10_cal = 16'b0000000001111000;
            15'd1344: log10_cal = 16'b0000000001111000;
            15'd1345: log10_cal = 16'b0000000001111001;
            15'd1346: log10_cal = 16'b0000000001111001;
            15'd1347: log10_cal = 16'b0000000001111001;
            15'd1348: log10_cal = 16'b0000000001111010;
            15'd1349: log10_cal = 16'b0000000001111010;
            15'd1350: log10_cal = 16'b0000000001111010;
            15'd1351: log10_cal = 16'b0000000001111011;
            15'd1352: log10_cal = 16'b0000000001111011;
            15'd1353: log10_cal = 16'b0000000001111011;
            15'd1354: log10_cal = 16'b0000000001111100;
            15'd1355: log10_cal = 16'b0000000001111100;
            15'd1356: log10_cal = 16'b0000000001111100;
            15'd1357: log10_cal = 16'b0000000001111101;
            15'd1358: log10_cal = 16'b0000000001111101;
            15'd1359: log10_cal = 16'b0000000001111101;
            15'd1360: log10_cal = 16'b0000000001111110;
            15'd1361: log10_cal = 16'b0000000001111110;
            15'd1362: log10_cal = 16'b0000000001111110;
            15'd1363: log10_cal = 16'b0000000001111111;
            15'd1364: log10_cal = 16'b0000000001111111;
            15'd1365: log10_cal = 16'b0000000001111111;
            15'd1366: log10_cal = 16'b0000000010000000;
            15'd1367: log10_cal = 16'b0000000010000000;
            15'd1368: log10_cal = 16'b0000000010000000;
            15'd1369: log10_cal = 16'b0000000010000001;
            15'd1370: log10_cal = 16'b0000000010000001;
            15'd1371: log10_cal = 16'b0000000010000001;
            15'd1372: log10_cal = 16'b0000000010000010;
            15'd1373: log10_cal = 16'b0000000010000010;
            15'd1374: log10_cal = 16'b0000000010000010;
            15'd1375: log10_cal = 16'b0000000010000011;
            15'd1376: log10_cal = 16'b0000000010000011;
            15'd1377: log10_cal = 16'b0000000010000011;
            15'd1378: log10_cal = 16'b0000000010000100;
            15'd1379: log10_cal = 16'b0000000010000100;
            15'd1380: log10_cal = 16'b0000000010000100;
            15'd1381: log10_cal = 16'b0000000010000101;
            15'd1382: log10_cal = 16'b0000000010000101;
            15'd1383: log10_cal = 16'b0000000010000101;
            15'd1384: log10_cal = 16'b0000000010000101;
            15'd1385: log10_cal = 16'b0000000010000110;
            15'd1386: log10_cal = 16'b0000000010000110;
            15'd1387: log10_cal = 16'b0000000010000110;
            15'd1388: log10_cal = 16'b0000000010000111;
            15'd1389: log10_cal = 16'b0000000010000111;
            15'd1390: log10_cal = 16'b0000000010000111;
            15'd1391: log10_cal = 16'b0000000010001000;
            15'd1392: log10_cal = 16'b0000000010001000;
            15'd1393: log10_cal = 16'b0000000010001000;
            15'd1394: log10_cal = 16'b0000000010001001;
            15'd1395: log10_cal = 16'b0000000010001001;
            15'd1396: log10_cal = 16'b0000000010001001;
            15'd1397: log10_cal = 16'b0000000010001010;
            15'd1398: log10_cal = 16'b0000000010001010;
            15'd1399: log10_cal = 16'b0000000010001010;
            15'd1400: log10_cal = 16'b0000000010001011;
            15'd1401: log10_cal = 16'b0000000010001011;
            15'd1402: log10_cal = 16'b0000000010001011;
            15'd1403: log10_cal = 16'b0000000010001100;
            15'd1404: log10_cal = 16'b0000000010001100;
            15'd1405: log10_cal = 16'b0000000010001100;
            15'd1406: log10_cal = 16'b0000000010001100;
            15'd1407: log10_cal = 16'b0000000010001101;
            15'd1408: log10_cal = 16'b0000000010001101;
            15'd1409: log10_cal = 16'b0000000010001101;
            15'd1410: log10_cal = 16'b0000000010001110;
            15'd1411: log10_cal = 16'b0000000010001110;
            15'd1412: log10_cal = 16'b0000000010001110;
            15'd1413: log10_cal = 16'b0000000010001111;
            15'd1414: log10_cal = 16'b0000000010001111;
            15'd1415: log10_cal = 16'b0000000010001111;
            15'd1416: log10_cal = 16'b0000000010010000;
            15'd1417: log10_cal = 16'b0000000010010000;
            15'd1418: log10_cal = 16'b0000000010010000;
            15'd1419: log10_cal = 16'b0000000010010001;
            15'd1420: log10_cal = 16'b0000000010010001;
            15'd1421: log10_cal = 16'b0000000010010001;
            15'd1422: log10_cal = 16'b0000000010010010;
            15'd1423: log10_cal = 16'b0000000010010010;
            15'd1424: log10_cal = 16'b0000000010010010;
            15'd1425: log10_cal = 16'b0000000010010010;
            15'd1426: log10_cal = 16'b0000000010010011;
            15'd1427: log10_cal = 16'b0000000010010011;
            15'd1428: log10_cal = 16'b0000000010010011;
            15'd1429: log10_cal = 16'b0000000010010100;
            15'd1430: log10_cal = 16'b0000000010010100;
            15'd1431: log10_cal = 16'b0000000010010100;
            15'd1432: log10_cal = 16'b0000000010010101;
            15'd1433: log10_cal = 16'b0000000010010101;
            15'd1434: log10_cal = 16'b0000000010010101;
            15'd1435: log10_cal = 16'b0000000010010110;
            15'd1436: log10_cal = 16'b0000000010010110;
            15'd1437: log10_cal = 16'b0000000010010110;
            15'd1438: log10_cal = 16'b0000000010010110;
            15'd1439: log10_cal = 16'b0000000010010111;
            15'd1440: log10_cal = 16'b0000000010010111;
            15'd1441: log10_cal = 16'b0000000010010111;
            15'd1442: log10_cal = 16'b0000000010011000;
            15'd1443: log10_cal = 16'b0000000010011000;
            15'd1444: log10_cal = 16'b0000000010011000;
            15'd1445: log10_cal = 16'b0000000010011001;
            15'd1446: log10_cal = 16'b0000000010011001;
            15'd1447: log10_cal = 16'b0000000010011001;
            15'd1448: log10_cal = 16'b0000000010011010;
            15'd1449: log10_cal = 16'b0000000010011010;
            15'd1450: log10_cal = 16'b0000000010011010;
            15'd1451: log10_cal = 16'b0000000010011011;
            15'd1452: log10_cal = 16'b0000000010011011;
            15'd1453: log10_cal = 16'b0000000010011011;
            15'd1454: log10_cal = 16'b0000000010011011;
            15'd1455: log10_cal = 16'b0000000010011100;
            15'd1456: log10_cal = 16'b0000000010011100;
            15'd1457: log10_cal = 16'b0000000010011100;
            15'd1458: log10_cal = 16'b0000000010011101;
            15'd1459: log10_cal = 16'b0000000010011101;
            15'd1460: log10_cal = 16'b0000000010011101;
            15'd1461: log10_cal = 16'b0000000010011110;
            15'd1462: log10_cal = 16'b0000000010011110;
            15'd1463: log10_cal = 16'b0000000010011110;
            15'd1464: log10_cal = 16'b0000000010011110;
            15'd1465: log10_cal = 16'b0000000010011111;
            15'd1466: log10_cal = 16'b0000000010011111;
            15'd1467: log10_cal = 16'b0000000010011111;
            15'd1468: log10_cal = 16'b0000000010100000;
            15'd1469: log10_cal = 16'b0000000010100000;
            15'd1470: log10_cal = 16'b0000000010100000;
            15'd1471: log10_cal = 16'b0000000010100001;
            15'd1472: log10_cal = 16'b0000000010100001;
            15'd1473: log10_cal = 16'b0000000010100001;
            15'd1474: log10_cal = 16'b0000000010100001;
            15'd1475: log10_cal = 16'b0000000010100010;
            15'd1476: log10_cal = 16'b0000000010100010;
            15'd1477: log10_cal = 16'b0000000010100010;
            15'd1478: log10_cal = 16'b0000000010100011;
            15'd1479: log10_cal = 16'b0000000010100011;
            15'd1480: log10_cal = 16'b0000000010100011;
            15'd1481: log10_cal = 16'b0000000010100100;
            15'd1482: log10_cal = 16'b0000000010100100;
            15'd1483: log10_cal = 16'b0000000010100100;
            15'd1484: log10_cal = 16'b0000000010100101;
            15'd1485: log10_cal = 16'b0000000010100101;
            15'd1486: log10_cal = 16'b0000000010100101;
            15'd1487: log10_cal = 16'b0000000010100101;
            15'd1488: log10_cal = 16'b0000000010100110;
            15'd1489: log10_cal = 16'b0000000010100110;
            15'd1490: log10_cal = 16'b0000000010100110;
            15'd1491: log10_cal = 16'b0000000010100111;
            15'd1492: log10_cal = 16'b0000000010100111;
            15'd1493: log10_cal = 16'b0000000010100111;
            15'd1494: log10_cal = 16'b0000000010100111;
            15'd1495: log10_cal = 16'b0000000010101000;
            15'd1496: log10_cal = 16'b0000000010101000;
            15'd1497: log10_cal = 16'b0000000010101000;
            15'd1498: log10_cal = 16'b0000000010101001;
            15'd1499: log10_cal = 16'b0000000010101001;
            15'd1500: log10_cal = 16'b0000000010101001;
            15'd1501: log10_cal = 16'b0000000010101010;
            15'd1502: log10_cal = 16'b0000000010101010;
            15'd1503: log10_cal = 16'b0000000010101010;
            15'd1504: log10_cal = 16'b0000000010101010;
            15'd1505: log10_cal = 16'b0000000010101011;
            15'd1506: log10_cal = 16'b0000000010101011;
            15'd1507: log10_cal = 16'b0000000010101011;
            15'd1508: log10_cal = 16'b0000000010101100;
            15'd1509: log10_cal = 16'b0000000010101100;
            15'd1510: log10_cal = 16'b0000000010101100;
            15'd1511: log10_cal = 16'b0000000010101101;
            15'd1512: log10_cal = 16'b0000000010101101;
            15'd1513: log10_cal = 16'b0000000010101101;
            15'd1514: log10_cal = 16'b0000000010101101;
            15'd1515: log10_cal = 16'b0000000010101110;
            15'd1516: log10_cal = 16'b0000000010101110;
            15'd1517: log10_cal = 16'b0000000010101110;
            15'd1518: log10_cal = 16'b0000000010101111;
            15'd1519: log10_cal = 16'b0000000010101111;
            15'd1520: log10_cal = 16'b0000000010101111;
            15'd1521: log10_cal = 16'b0000000010101111;
            15'd1522: log10_cal = 16'b0000000010110000;
            15'd1523: log10_cal = 16'b0000000010110000;
            15'd1524: log10_cal = 16'b0000000010110000;
            15'd1525: log10_cal = 16'b0000000010110001;
            15'd1526: log10_cal = 16'b0000000010110001;
            15'd1527: log10_cal = 16'b0000000010110001;
            15'd1528: log10_cal = 16'b0000000010110001;
            15'd1529: log10_cal = 16'b0000000010110010;
            15'd1530: log10_cal = 16'b0000000010110010;
            15'd1531: log10_cal = 16'b0000000010110010;
            15'd1532: log10_cal = 16'b0000000010110011;
            15'd1533: log10_cal = 16'b0000000010110011;
            15'd1534: log10_cal = 16'b0000000010110011;
            15'd1535: log10_cal = 16'b0000000010110100;
            15'd1536: log10_cal = 16'b0000000010110100;
            15'd1537: log10_cal = 16'b0000000010110100;
            15'd1538: log10_cal = 16'b0000000010110100;
            15'd1539: log10_cal = 16'b0000000010110101;
            15'd1540: log10_cal = 16'b0000000010110101;
            15'd1541: log10_cal = 16'b0000000010110101;
            15'd1542: log10_cal = 16'b0000000010110110;
            15'd1543: log10_cal = 16'b0000000010110110;
            15'd1544: log10_cal = 16'b0000000010110110;
            15'd1545: log10_cal = 16'b0000000010110110;
            15'd1546: log10_cal = 16'b0000000010110111;
            15'd1547: log10_cal = 16'b0000000010110111;
            15'd1548: log10_cal = 16'b0000000010110111;
            15'd1549: log10_cal = 16'b0000000010111000;
            15'd1550: log10_cal = 16'b0000000010111000;
            15'd1551: log10_cal = 16'b0000000010111000;
            15'd1552: log10_cal = 16'b0000000010111000;
            15'd1553: log10_cal = 16'b0000000010111001;
            15'd1554: log10_cal = 16'b0000000010111001;
            15'd1555: log10_cal = 16'b0000000010111001;
            15'd1556: log10_cal = 16'b0000000010111010;
            15'd1557: log10_cal = 16'b0000000010111010;
            15'd1558: log10_cal = 16'b0000000010111010;
            15'd1559: log10_cal = 16'b0000000010111010;
            15'd1560: log10_cal = 16'b0000000010111011;
            15'd1561: log10_cal = 16'b0000000010111011;
            15'd1562: log10_cal = 16'b0000000010111011;
            15'd1563: log10_cal = 16'b0000000010111100;
            15'd1564: log10_cal = 16'b0000000010111100;
            15'd1565: log10_cal = 16'b0000000010111100;
            15'd1566: log10_cal = 16'b0000000010111100;
            15'd1567: log10_cal = 16'b0000000010111101;
            15'd1568: log10_cal = 16'b0000000010111101;
            15'd1569: log10_cal = 16'b0000000010111101;
            15'd1570: log10_cal = 16'b0000000010111110;
            15'd1571: log10_cal = 16'b0000000010111110;
            15'd1572: log10_cal = 16'b0000000010111110;
            15'd1573: log10_cal = 16'b0000000010111110;
            15'd1574: log10_cal = 16'b0000000010111111;
            15'd1575: log10_cal = 16'b0000000010111111;
            15'd1576: log10_cal = 16'b0000000010111111;
            15'd1577: log10_cal = 16'b0000000011000000;
            15'd1578: log10_cal = 16'b0000000011000000;
            15'd1579: log10_cal = 16'b0000000011000000;
            15'd1580: log10_cal = 16'b0000000011000000;
            15'd1581: log10_cal = 16'b0000000011000001;
            15'd1582: log10_cal = 16'b0000000011000001;
            15'd1583: log10_cal = 16'b0000000011000001;
            15'd1584: log10_cal = 16'b0000000011000010;
            15'd1585: log10_cal = 16'b0000000011000010;
            15'd1586: log10_cal = 16'b0000000011000010;
            15'd1587: log10_cal = 16'b0000000011000010;
            15'd1588: log10_cal = 16'b0000000011000011;
            15'd1589: log10_cal = 16'b0000000011000011;
            15'd1590: log10_cal = 16'b0000000011000011;
            15'd1591: log10_cal = 16'b0000000011000011;
            15'd1592: log10_cal = 16'b0000000011000100;
            15'd1593: log10_cal = 16'b0000000011000100;
            15'd1594: log10_cal = 16'b0000000011000100;
            15'd1595: log10_cal = 16'b0000000011000101;
            15'd1596: log10_cal = 16'b0000000011000101;
            15'd1597: log10_cal = 16'b0000000011000101;
            15'd1598: log10_cal = 16'b0000000011000101;
            15'd1599: log10_cal = 16'b0000000011000110;
            15'd1600: log10_cal = 16'b0000000011000110;
            15'd1601: log10_cal = 16'b0000000011000110;
            15'd1602: log10_cal = 16'b0000000011000111;
            15'd1603: log10_cal = 16'b0000000011000111;
            15'd1604: log10_cal = 16'b0000000011000111;
            15'd1605: log10_cal = 16'b0000000011000111;
            15'd1606: log10_cal = 16'b0000000011001000;
            15'd1607: log10_cal = 16'b0000000011001000;
            15'd1608: log10_cal = 16'b0000000011001000;
            15'd1609: log10_cal = 16'b0000000011001000;
            15'd1610: log10_cal = 16'b0000000011001001;
            15'd1611: log10_cal = 16'b0000000011001001;
            15'd1612: log10_cal = 16'b0000000011001001;
            15'd1613: log10_cal = 16'b0000000011001010;
            15'd1614: log10_cal = 16'b0000000011001010;
            15'd1615: log10_cal = 16'b0000000011001010;
            15'd1616: log10_cal = 16'b0000000011001010;
            15'd1617: log10_cal = 16'b0000000011001011;
            15'd1618: log10_cal = 16'b0000000011001011;
            15'd1619: log10_cal = 16'b0000000011001011;
            15'd1620: log10_cal = 16'b0000000011001011;
            15'd1621: log10_cal = 16'b0000000011001100;
            15'd1622: log10_cal = 16'b0000000011001100;
            15'd1623: log10_cal = 16'b0000000011001100;
            15'd1624: log10_cal = 16'b0000000011001101;
            15'd1625: log10_cal = 16'b0000000011001101;
            15'd1626: log10_cal = 16'b0000000011001101;
            15'd1627: log10_cal = 16'b0000000011001101;
            15'd1628: log10_cal = 16'b0000000011001110;
            15'd1629: log10_cal = 16'b0000000011001110;
            15'd1630: log10_cal = 16'b0000000011001110;
            15'd1631: log10_cal = 16'b0000000011001111;
            15'd1632: log10_cal = 16'b0000000011001111;
            15'd1633: log10_cal = 16'b0000000011001111;
            15'd1634: log10_cal = 16'b0000000011001111;
            15'd1635: log10_cal = 16'b0000000011010000;
            15'd1636: log10_cal = 16'b0000000011010000;
            15'd1637: log10_cal = 16'b0000000011010000;
            15'd1638: log10_cal = 16'b0000000011010000;
            15'd1639: log10_cal = 16'b0000000011010001;
            15'd1640: log10_cal = 16'b0000000011010001;
            15'd1641: log10_cal = 16'b0000000011010001;
            15'd1642: log10_cal = 16'b0000000011010001;
            15'd1643: log10_cal = 16'b0000000011010010;
            15'd1644: log10_cal = 16'b0000000011010010;
            15'd1645: log10_cal = 16'b0000000011010010;
            15'd1646: log10_cal = 16'b0000000011010011;
            15'd1647: log10_cal = 16'b0000000011010011;
            15'd1648: log10_cal = 16'b0000000011010011;
            15'd1649: log10_cal = 16'b0000000011010011;
            15'd1650: log10_cal = 16'b0000000011010100;
            15'd1651: log10_cal = 16'b0000000011010100;
            15'd1652: log10_cal = 16'b0000000011010100;
            15'd1653: log10_cal = 16'b0000000011010100;
            15'd1654: log10_cal = 16'b0000000011010101;
            15'd1655: log10_cal = 16'b0000000011010101;
            15'd1656: log10_cal = 16'b0000000011010101;
            15'd1657: log10_cal = 16'b0000000011010110;
            15'd1658: log10_cal = 16'b0000000011010110;
            15'd1659: log10_cal = 16'b0000000011010110;
            15'd1660: log10_cal = 16'b0000000011010110;
            15'd1661: log10_cal = 16'b0000000011010111;
            15'd1662: log10_cal = 16'b0000000011010111;
            15'd1663: log10_cal = 16'b0000000011010111;
            15'd1664: log10_cal = 16'b0000000011010111;
            15'd1665: log10_cal = 16'b0000000011011000;
            15'd1666: log10_cal = 16'b0000000011011000;
            15'd1667: log10_cal = 16'b0000000011011000;
            15'd1668: log10_cal = 16'b0000000011011000;
            15'd1669: log10_cal = 16'b0000000011011001;
            15'd1670: log10_cal = 16'b0000000011011001;
            15'd1671: log10_cal = 16'b0000000011011001;
            15'd1672: log10_cal = 16'b0000000011011010;
            15'd1673: log10_cal = 16'b0000000011011010;
            15'd1674: log10_cal = 16'b0000000011011010;
            15'd1675: log10_cal = 16'b0000000011011010;
            15'd1676: log10_cal = 16'b0000000011011011;
            15'd1677: log10_cal = 16'b0000000011011011;
            15'd1678: log10_cal = 16'b0000000011011011;
            15'd1679: log10_cal = 16'b0000000011011011;
            15'd1680: log10_cal = 16'b0000000011011100;
            15'd1681: log10_cal = 16'b0000000011011100;
            15'd1682: log10_cal = 16'b0000000011011100;
            15'd1683: log10_cal = 16'b0000000011011100;
            15'd1684: log10_cal = 16'b0000000011011101;
            15'd1685: log10_cal = 16'b0000000011011101;
            15'd1686: log10_cal = 16'b0000000011011101;
            15'd1687: log10_cal = 16'b0000000011011110;
            15'd1688: log10_cal = 16'b0000000011011110;
            15'd1689: log10_cal = 16'b0000000011011110;
            15'd1690: log10_cal = 16'b0000000011011110;
            15'd1691: log10_cal = 16'b0000000011011111;
            15'd1692: log10_cal = 16'b0000000011011111;
            15'd1693: log10_cal = 16'b0000000011011111;
            15'd1694: log10_cal = 16'b0000000011011111;
            15'd1695: log10_cal = 16'b0000000011100000;
            15'd1696: log10_cal = 16'b0000000011100000;
            15'd1697: log10_cal = 16'b0000000011100000;
            15'd1698: log10_cal = 16'b0000000011100000;
            15'd1699: log10_cal = 16'b0000000011100001;
            15'd1700: log10_cal = 16'b0000000011100001;
            15'd1701: log10_cal = 16'b0000000011100001;
            15'd1702: log10_cal = 16'b0000000011100001;
            15'd1703: log10_cal = 16'b0000000011100010;
            15'd1704: log10_cal = 16'b0000000011100010;
            15'd1705: log10_cal = 16'b0000000011100010;
            15'd1706: log10_cal = 16'b0000000011100010;
            15'd1707: log10_cal = 16'b0000000011100011;
            15'd1708: log10_cal = 16'b0000000011100011;
            15'd1709: log10_cal = 16'b0000000011100011;
            15'd1710: log10_cal = 16'b0000000011100100;
            15'd1711: log10_cal = 16'b0000000011100100;
            15'd1712: log10_cal = 16'b0000000011100100;
            15'd1713: log10_cal = 16'b0000000011100100;
            15'd1714: log10_cal = 16'b0000000011100101;
            15'd1715: log10_cal = 16'b0000000011100101;
            15'd1716: log10_cal = 16'b0000000011100101;
            15'd1717: log10_cal = 16'b0000000011100101;
            15'd1718: log10_cal = 16'b0000000011100110;
            15'd1719: log10_cal = 16'b0000000011100110;
            15'd1720: log10_cal = 16'b0000000011100110;
            15'd1721: log10_cal = 16'b0000000011100110;
            15'd1722: log10_cal = 16'b0000000011100111;
            15'd1723: log10_cal = 16'b0000000011100111;
            15'd1724: log10_cal = 16'b0000000011100111;
            15'd1725: log10_cal = 16'b0000000011100111;
            15'd1726: log10_cal = 16'b0000000011101000;
            15'd1727: log10_cal = 16'b0000000011101000;
            15'd1728: log10_cal = 16'b0000000011101000;
            15'd1729: log10_cal = 16'b0000000011101000;
            15'd1730: log10_cal = 16'b0000000011101001;
            15'd1731: log10_cal = 16'b0000000011101001;
            15'd1732: log10_cal = 16'b0000000011101001;
            15'd1733: log10_cal = 16'b0000000011101001;
            15'd1734: log10_cal = 16'b0000000011101010;
            15'd1735: log10_cal = 16'b0000000011101010;
            15'd1736: log10_cal = 16'b0000000011101010;
            15'd1737: log10_cal = 16'b0000000011101011;
            15'd1738: log10_cal = 16'b0000000011101011;
            15'd1739: log10_cal = 16'b0000000011101011;
            15'd1740: log10_cal = 16'b0000000011101011;
            15'd1741: log10_cal = 16'b0000000011101100;
            15'd1742: log10_cal = 16'b0000000011101100;
            15'd1743: log10_cal = 16'b0000000011101100;
            15'd1744: log10_cal = 16'b0000000011101100;
            15'd1745: log10_cal = 16'b0000000011101101;
            15'd1746: log10_cal = 16'b0000000011101101;
            15'd1747: log10_cal = 16'b0000000011101101;
            15'd1748: log10_cal = 16'b0000000011101101;
            15'd1749: log10_cal = 16'b0000000011101110;
            15'd1750: log10_cal = 16'b0000000011101110;
            15'd1751: log10_cal = 16'b0000000011101110;
            15'd1752: log10_cal = 16'b0000000011101110;
            15'd1753: log10_cal = 16'b0000000011101111;
            15'd1754: log10_cal = 16'b0000000011101111;
            15'd1755: log10_cal = 16'b0000000011101111;
            15'd1756: log10_cal = 16'b0000000011101111;
            15'd1757: log10_cal = 16'b0000000011110000;
            15'd1758: log10_cal = 16'b0000000011110000;
            15'd1759: log10_cal = 16'b0000000011110000;
            15'd1760: log10_cal = 16'b0000000011110000;
            15'd1761: log10_cal = 16'b0000000011110001;
            15'd1762: log10_cal = 16'b0000000011110001;
            15'd1763: log10_cal = 16'b0000000011110001;
            15'd1764: log10_cal = 16'b0000000011110001;
            15'd1765: log10_cal = 16'b0000000011110010;
            15'd1766: log10_cal = 16'b0000000011110010;
            15'd1767: log10_cal = 16'b0000000011110010;
            15'd1768: log10_cal = 16'b0000000011110010;
            15'd1769: log10_cal = 16'b0000000011110011;
            15'd1770: log10_cal = 16'b0000000011110011;
            15'd1771: log10_cal = 16'b0000000011110011;
            15'd1772: log10_cal = 16'b0000000011110011;
            15'd1773: log10_cal = 16'b0000000011110100;
            15'd1774: log10_cal = 16'b0000000011110100;
            15'd1775: log10_cal = 16'b0000000011110100;
            15'd1776: log10_cal = 16'b0000000011110100;
            15'd1777: log10_cal = 16'b0000000011110101;
            15'd1778: log10_cal = 16'b0000000011110101;
            15'd1779: log10_cal = 16'b0000000011110101;
            15'd1780: log10_cal = 16'b0000000011110101;
            15'd1781: log10_cal = 16'b0000000011110110;
            15'd1782: log10_cal = 16'b0000000011110110;
            15'd1783: log10_cal = 16'b0000000011110110;
            15'd1784: log10_cal = 16'b0000000011110110;
            15'd1785: log10_cal = 16'b0000000011110111;
            15'd1786: log10_cal = 16'b0000000011110111;
            15'd1787: log10_cal = 16'b0000000011110111;
            15'd1788: log10_cal = 16'b0000000011110111;
            15'd1789: log10_cal = 16'b0000000011111000;
            15'd1790: log10_cal = 16'b0000000011111000;
            15'd1791: log10_cal = 16'b0000000011111000;
            15'd1792: log10_cal = 16'b0000000011111000;
            15'd1793: log10_cal = 16'b0000000011111001;
            15'd1794: log10_cal = 16'b0000000011111001;
            15'd1795: log10_cal = 16'b0000000011111001;
            15'd1796: log10_cal = 16'b0000000011111001;
            15'd1797: log10_cal = 16'b0000000011111010;
            15'd1798: log10_cal = 16'b0000000011111010;
            15'd1799: log10_cal = 16'b0000000011111010;
            15'd1800: log10_cal = 16'b0000000011111010;
            15'd1801: log10_cal = 16'b0000000011111011;
            15'd1802: log10_cal = 16'b0000000011111011;
            15'd1803: log10_cal = 16'b0000000011111011;
            15'd1804: log10_cal = 16'b0000000011111011;
            15'd1805: log10_cal = 16'b0000000011111100;
            15'd1806: log10_cal = 16'b0000000011111100;
            15'd1807: log10_cal = 16'b0000000011111100;
            15'd1808: log10_cal = 16'b0000000011111100;
            15'd1809: log10_cal = 16'b0000000011111101;
            15'd1810: log10_cal = 16'b0000000011111101;
            15'd1811: log10_cal = 16'b0000000011111101;
            15'd1812: log10_cal = 16'b0000000011111101;
            15'd1813: log10_cal = 16'b0000000011111110;
            15'd1814: log10_cal = 16'b0000000011111110;
            15'd1815: log10_cal = 16'b0000000011111110;
            15'd1816: log10_cal = 16'b0000000011111110;
            15'd1817: log10_cal = 16'b0000000011111111;
            15'd1818: log10_cal = 16'b0000000011111111;
            15'd1819: log10_cal = 16'b0000000011111111;
            15'd1820: log10_cal = 16'b0000000011111111;
            15'd1821: log10_cal = 16'b0000000100000000;
            15'd1822: log10_cal = 16'b0000000100000000;
            15'd1823: log10_cal = 16'b0000000100000000;
            15'd1824: log10_cal = 16'b0000000100000000;
            15'd1825: log10_cal = 16'b0000000100000000;
            15'd1826: log10_cal = 16'b0000000100000001;
            15'd1827: log10_cal = 16'b0000000100000001;
            15'd1828: log10_cal = 16'b0000000100000001;
            15'd1829: log10_cal = 16'b0000000100000001;
            15'd1830: log10_cal = 16'b0000000100000010;
            15'd1831: log10_cal = 16'b0000000100000010;
            15'd1832: log10_cal = 16'b0000000100000010;
            15'd1833: log10_cal = 16'b0000000100000010;
            15'd1834: log10_cal = 16'b0000000100000011;
            15'd1835: log10_cal = 16'b0000000100000011;
            15'd1836: log10_cal = 16'b0000000100000011;
            15'd1837: log10_cal = 16'b0000000100000011;
            15'd1838: log10_cal = 16'b0000000100000100;
            15'd1839: log10_cal = 16'b0000000100000100;
            15'd1840: log10_cal = 16'b0000000100000100;
            15'd1841: log10_cal = 16'b0000000100000100;
            15'd1842: log10_cal = 16'b0000000100000101;
            15'd1843: log10_cal = 16'b0000000100000101;
            15'd1844: log10_cal = 16'b0000000100000101;
            15'd1845: log10_cal = 16'b0000000100000101;
            15'd1846: log10_cal = 16'b0000000100000110;
            15'd1847: log10_cal = 16'b0000000100000110;
            15'd1848: log10_cal = 16'b0000000100000110;
            15'd1849: log10_cal = 16'b0000000100000110;
            15'd1850: log10_cal = 16'b0000000100000111;
            15'd1851: log10_cal = 16'b0000000100000111;
            15'd1852: log10_cal = 16'b0000000100000111;
            15'd1853: log10_cal = 16'b0000000100000111;
            15'd1854: log10_cal = 16'b0000000100000111;
            15'd1855: log10_cal = 16'b0000000100001000;
            15'd1856: log10_cal = 16'b0000000100001000;
            15'd1857: log10_cal = 16'b0000000100001000;
            15'd1858: log10_cal = 16'b0000000100001000;
            15'd1859: log10_cal = 16'b0000000100001001;
            15'd1860: log10_cal = 16'b0000000100001001;
            15'd1861: log10_cal = 16'b0000000100001001;
            15'd1862: log10_cal = 16'b0000000100001001;
            15'd1863: log10_cal = 16'b0000000100001010;
            15'd1864: log10_cal = 16'b0000000100001010;
            15'd1865: log10_cal = 16'b0000000100001010;
            15'd1866: log10_cal = 16'b0000000100001010;
            15'd1867: log10_cal = 16'b0000000100001011;
            15'd1868: log10_cal = 16'b0000000100001011;
            15'd1869: log10_cal = 16'b0000000100001011;
            15'd1870: log10_cal = 16'b0000000100001011;
            15'd1871: log10_cal = 16'b0000000100001100;
            15'd1872: log10_cal = 16'b0000000100001100;
            15'd1873: log10_cal = 16'b0000000100001100;
            15'd1874: log10_cal = 16'b0000000100001100;
            15'd1875: log10_cal = 16'b0000000100001101;
            15'd1876: log10_cal = 16'b0000000100001101;
            15'd1877: log10_cal = 16'b0000000100001101;
            15'd1878: log10_cal = 16'b0000000100001101;
            15'd1879: log10_cal = 16'b0000000100001101;
            15'd1880: log10_cal = 16'b0000000100001110;
            15'd1881: log10_cal = 16'b0000000100001110;
            15'd1882: log10_cal = 16'b0000000100001110;
            15'd1883: log10_cal = 16'b0000000100001110;
            15'd1884: log10_cal = 16'b0000000100001111;
            15'd1885: log10_cal = 16'b0000000100001111;
            15'd1886: log10_cal = 16'b0000000100001111;
            15'd1887: log10_cal = 16'b0000000100001111;
            15'd1888: log10_cal = 16'b0000000100010000;
            15'd1889: log10_cal = 16'b0000000100010000;
            15'd1890: log10_cal = 16'b0000000100010000;
            15'd1891: log10_cal = 16'b0000000100010000;
            15'd1892: log10_cal = 16'b0000000100010001;
            15'd1893: log10_cal = 16'b0000000100010001;
            15'd1894: log10_cal = 16'b0000000100010001;
            15'd1895: log10_cal = 16'b0000000100010001;
            15'd1896: log10_cal = 16'b0000000100010001;
            15'd1897: log10_cal = 16'b0000000100010010;
            15'd1898: log10_cal = 16'b0000000100010010;
            15'd1899: log10_cal = 16'b0000000100010010;
            15'd1900: log10_cal = 16'b0000000100010010;
            15'd1901: log10_cal = 16'b0000000100010011;
            15'd1902: log10_cal = 16'b0000000100010011;
            15'd1903: log10_cal = 16'b0000000100010011;
            15'd1904: log10_cal = 16'b0000000100010011;
            15'd1905: log10_cal = 16'b0000000100010100;
            15'd1906: log10_cal = 16'b0000000100010100;
            15'd1907: log10_cal = 16'b0000000100010100;
            15'd1908: log10_cal = 16'b0000000100010100;
            15'd1909: log10_cal = 16'b0000000100010100;
            15'd1910: log10_cal = 16'b0000000100010101;
            15'd1911: log10_cal = 16'b0000000100010101;
            15'd1912: log10_cal = 16'b0000000100010101;
            15'd1913: log10_cal = 16'b0000000100010101;
            15'd1914: log10_cal = 16'b0000000100010110;
            15'd1915: log10_cal = 16'b0000000100010110;
            15'd1916: log10_cal = 16'b0000000100010110;
            15'd1917: log10_cal = 16'b0000000100010110;
            15'd1918: log10_cal = 16'b0000000100010111;
            15'd1919: log10_cal = 16'b0000000100010111;
            15'd1920: log10_cal = 16'b0000000100010111;
            15'd1921: log10_cal = 16'b0000000100010111;
            15'd1922: log10_cal = 16'b0000000100011000;
            15'd1923: log10_cal = 16'b0000000100011000;
            15'd1924: log10_cal = 16'b0000000100011000;
            15'd1925: log10_cal = 16'b0000000100011000;
            15'd1926: log10_cal = 16'b0000000100011000;
            15'd1927: log10_cal = 16'b0000000100011001;
            15'd1928: log10_cal = 16'b0000000100011001;
            15'd1929: log10_cal = 16'b0000000100011001;
            15'd1930: log10_cal = 16'b0000000100011001;
            15'd1931: log10_cal = 16'b0000000100011010;
            15'd1932: log10_cal = 16'b0000000100011010;
            15'd1933: log10_cal = 16'b0000000100011010;
            15'd1934: log10_cal = 16'b0000000100011010;
            15'd1935: log10_cal = 16'b0000000100011011;
            15'd1936: log10_cal = 16'b0000000100011011;
            15'd1937: log10_cal = 16'b0000000100011011;
            15'd1938: log10_cal = 16'b0000000100011011;
            15'd1939: log10_cal = 16'b0000000100011011;
            15'd1940: log10_cal = 16'b0000000100011100;
            15'd1941: log10_cal = 16'b0000000100011100;
            15'd1942: log10_cal = 16'b0000000100011100;
            15'd1943: log10_cal = 16'b0000000100011100;
            15'd1944: log10_cal = 16'b0000000100011101;
            15'd1945: log10_cal = 16'b0000000100011101;
            15'd1946: log10_cal = 16'b0000000100011101;
            15'd1947: log10_cal = 16'b0000000100011101;
            15'd1948: log10_cal = 16'b0000000100011101;
            15'd1949: log10_cal = 16'b0000000100011110;
            15'd1950: log10_cal = 16'b0000000100011110;
            15'd1951: log10_cal = 16'b0000000100011110;
            15'd1952: log10_cal = 16'b0000000100011110;
            15'd1953: log10_cal = 16'b0000000100011111;
            15'd1954: log10_cal = 16'b0000000100011111;
            15'd1955: log10_cal = 16'b0000000100011111;
            15'd1956: log10_cal = 16'b0000000100011111;
            15'd1957: log10_cal = 16'b0000000100100000;
            15'd1958: log10_cal = 16'b0000000100100000;
            15'd1959: log10_cal = 16'b0000000100100000;
            15'd1960: log10_cal = 16'b0000000100100000;
            15'd1961: log10_cal = 16'b0000000100100000;
            15'd1962: log10_cal = 16'b0000000100100001;
            15'd1963: log10_cal = 16'b0000000100100001;
            15'd1964: log10_cal = 16'b0000000100100001;
            15'd1965: log10_cal = 16'b0000000100100001;
            15'd1966: log10_cal = 16'b0000000100100010;
            15'd1967: log10_cal = 16'b0000000100100010;
            15'd1968: log10_cal = 16'b0000000100100010;
            15'd1969: log10_cal = 16'b0000000100100010;
            15'd1970: log10_cal = 16'b0000000100100010;
            15'd1971: log10_cal = 16'b0000000100100011;
            15'd1972: log10_cal = 16'b0000000100100011;
            15'd1973: log10_cal = 16'b0000000100100011;
            15'd1974: log10_cal = 16'b0000000100100011;
            15'd1975: log10_cal = 16'b0000000100100100;
            15'd1976: log10_cal = 16'b0000000100100100;
            15'd1977: log10_cal = 16'b0000000100100100;
            15'd1978: log10_cal = 16'b0000000100100100;
            15'd1979: log10_cal = 16'b0000000100100101;
            15'd1980: log10_cal = 16'b0000000100100101;
            15'd1981: log10_cal = 16'b0000000100100101;
            15'd1982: log10_cal = 16'b0000000100100101;
            15'd1983: log10_cal = 16'b0000000100100101;
            15'd1984: log10_cal = 16'b0000000100100110;
            15'd1985: log10_cal = 16'b0000000100100110;
            15'd1986: log10_cal = 16'b0000000100100110;
            15'd1987: log10_cal = 16'b0000000100100110;
            15'd1988: log10_cal = 16'b0000000100100111;
            15'd1989: log10_cal = 16'b0000000100100111;
            15'd1990: log10_cal = 16'b0000000100100111;
            15'd1991: log10_cal = 16'b0000000100100111;
            15'd1992: log10_cal = 16'b0000000100100111;
            15'd1993: log10_cal = 16'b0000000100101000;
            15'd1994: log10_cal = 16'b0000000100101000;
            15'd1995: log10_cal = 16'b0000000100101000;
            15'd1996: log10_cal = 16'b0000000100101000;
            15'd1997: log10_cal = 16'b0000000100101001;
            15'd1998: log10_cal = 16'b0000000100101001;
            15'd1999: log10_cal = 16'b0000000100101001;
            15'd2000: log10_cal = 16'b0000000100101001;
            15'd2001: log10_cal = 16'b0000000100101001;
            15'd2002: log10_cal = 16'b0000000100101010;
            15'd2003: log10_cal = 16'b0000000100101010;
            15'd2004: log10_cal = 16'b0000000100101010;
            15'd2005: log10_cal = 16'b0000000100101010;
            15'd2006: log10_cal = 16'b0000000100101011;
            15'd2007: log10_cal = 16'b0000000100101011;
            15'd2008: log10_cal = 16'b0000000100101011;
            15'd2009: log10_cal = 16'b0000000100101011;
            15'd2010: log10_cal = 16'b0000000100101011;
            15'd2011: log10_cal = 16'b0000000100101100;
            15'd2012: log10_cal = 16'b0000000100101100;
            15'd2013: log10_cal = 16'b0000000100101100;
            15'd2014: log10_cal = 16'b0000000100101100;
            15'd2015: log10_cal = 16'b0000000100101101;
            15'd2016: log10_cal = 16'b0000000100101101;
            15'd2017: log10_cal = 16'b0000000100101101;
            15'd2018: log10_cal = 16'b0000000100101101;
            15'd2019: log10_cal = 16'b0000000100101101;
            15'd2020: log10_cal = 16'b0000000100101110;
            15'd2021: log10_cal = 16'b0000000100101110;
            15'd2022: log10_cal = 16'b0000000100101110;
            15'd2023: log10_cal = 16'b0000000100101110;
            15'd2024: log10_cal = 16'b0000000100101111;
            15'd2025: log10_cal = 16'b0000000100101111;
            15'd2026: log10_cal = 16'b0000000100101111;
            15'd2027: log10_cal = 16'b0000000100101111;
            15'd2028: log10_cal = 16'b0000000100101111;
            15'd2029: log10_cal = 16'b0000000100110000;
            15'd2030: log10_cal = 16'b0000000100110000;
            15'd2031: log10_cal = 16'b0000000100110000;
            15'd2032: log10_cal = 16'b0000000100110000;
            15'd2033: log10_cal = 16'b0000000100110000;
            15'd2034: log10_cal = 16'b0000000100110001;
            15'd2035: log10_cal = 16'b0000000100110001;
            15'd2036: log10_cal = 16'b0000000100110001;
            15'd2037: log10_cal = 16'b0000000100110001;
            15'd2038: log10_cal = 16'b0000000100110010;
            15'd2039: log10_cal = 16'b0000000100110010;
            15'd2040: log10_cal = 16'b0000000100110010;
            15'd2041: log10_cal = 16'b0000000100110010;
            15'd2042: log10_cal = 16'b0000000100110010;
            15'd2043: log10_cal = 16'b0000000100110011;
            15'd2044: log10_cal = 16'b0000000100110011;
            15'd2045: log10_cal = 16'b0000000100110011;
            15'd2046: log10_cal = 16'b0000000100110011;
            15'd2047: log10_cal = 16'b0000000100110100;
            15'd2048: log10_cal = 16'b0000000100110100;
            15'd2049: log10_cal = 16'b0000000100110100;
            15'd2050: log10_cal = 16'b0000000100110100;
            15'd2051: log10_cal = 16'b0000000100110100;
            15'd2052: log10_cal = 16'b0000000100110101;
            15'd2053: log10_cal = 16'b0000000100110101;
            15'd2054: log10_cal = 16'b0000000100110101;
            15'd2055: log10_cal = 16'b0000000100110101;
            15'd2056: log10_cal = 16'b0000000100110101;
            15'd2057: log10_cal = 16'b0000000100110110;
            15'd2058: log10_cal = 16'b0000000100110110;
            15'd2059: log10_cal = 16'b0000000100110110;
            15'd2060: log10_cal = 16'b0000000100110110;
            15'd2061: log10_cal = 16'b0000000100110111;
            15'd2062: log10_cal = 16'b0000000100110111;
            15'd2063: log10_cal = 16'b0000000100110111;
            15'd2064: log10_cal = 16'b0000000100110111;
            15'd2065: log10_cal = 16'b0000000100110111;
            15'd2066: log10_cal = 16'b0000000100111000;
            15'd2067: log10_cal = 16'b0000000100111000;
            15'd2068: log10_cal = 16'b0000000100111000;
            15'd2069: log10_cal = 16'b0000000100111000;
            15'd2070: log10_cal = 16'b0000000100111001;
            15'd2071: log10_cal = 16'b0000000100111001;
            15'd2072: log10_cal = 16'b0000000100111001;
            15'd2073: log10_cal = 16'b0000000100111001;
            15'd2074: log10_cal = 16'b0000000100111001;
            15'd2075: log10_cal = 16'b0000000100111010;
            15'd2076: log10_cal = 16'b0000000100111010;
            15'd2077: log10_cal = 16'b0000000100111010;
            15'd2078: log10_cal = 16'b0000000100111010;
            15'd2079: log10_cal = 16'b0000000100111010;
            15'd2080: log10_cal = 16'b0000000100111011;
            15'd2081: log10_cal = 16'b0000000100111011;
            15'd2082: log10_cal = 16'b0000000100111011;
            15'd2083: log10_cal = 16'b0000000100111011;
            15'd2084: log10_cal = 16'b0000000100111100;
            15'd2085: log10_cal = 16'b0000000100111100;
            15'd2086: log10_cal = 16'b0000000100111100;
            15'd2087: log10_cal = 16'b0000000100111100;
            15'd2088: log10_cal = 16'b0000000100111100;
            15'd2089: log10_cal = 16'b0000000100111101;
            15'd2090: log10_cal = 16'b0000000100111101;
            15'd2091: log10_cal = 16'b0000000100111101;
            15'd2092: log10_cal = 16'b0000000100111101;
            15'd2093: log10_cal = 16'b0000000100111101;
            15'd2094: log10_cal = 16'b0000000100111110;
            15'd2095: log10_cal = 16'b0000000100111110;
            15'd2096: log10_cal = 16'b0000000100111110;
            15'd2097: log10_cal = 16'b0000000100111110;
            15'd2098: log10_cal = 16'b0000000100111110;
            15'd2099: log10_cal = 16'b0000000100111111;
            15'd2100: log10_cal = 16'b0000000100111111;
            15'd2101: log10_cal = 16'b0000000100111111;
            15'd2102: log10_cal = 16'b0000000100111111;
            15'd2103: log10_cal = 16'b0000000101000000;
            15'd2104: log10_cal = 16'b0000000101000000;
            15'd2105: log10_cal = 16'b0000000101000000;
            15'd2106: log10_cal = 16'b0000000101000000;
            15'd2107: log10_cal = 16'b0000000101000000;
            15'd2108: log10_cal = 16'b0000000101000001;
            15'd2109: log10_cal = 16'b0000000101000001;
            15'd2110: log10_cal = 16'b0000000101000001;
            15'd2111: log10_cal = 16'b0000000101000001;
            15'd2112: log10_cal = 16'b0000000101000001;
            15'd2113: log10_cal = 16'b0000000101000010;
            15'd2114: log10_cal = 16'b0000000101000010;
            15'd2115: log10_cal = 16'b0000000101000010;
            15'd2116: log10_cal = 16'b0000000101000010;
            15'd2117: log10_cal = 16'b0000000101000010;
            15'd2118: log10_cal = 16'b0000000101000011;
            15'd2119: log10_cal = 16'b0000000101000011;
            15'd2120: log10_cal = 16'b0000000101000011;
            15'd2121: log10_cal = 16'b0000000101000011;
            15'd2122: log10_cal = 16'b0000000101000100;
            15'd2123: log10_cal = 16'b0000000101000100;
            15'd2124: log10_cal = 16'b0000000101000100;
            15'd2125: log10_cal = 16'b0000000101000100;
            15'd2126: log10_cal = 16'b0000000101000100;
            15'd2127: log10_cal = 16'b0000000101000101;
            15'd2128: log10_cal = 16'b0000000101000101;
            15'd2129: log10_cal = 16'b0000000101000101;
            15'd2130: log10_cal = 16'b0000000101000101;
            15'd2131: log10_cal = 16'b0000000101000101;
            15'd2132: log10_cal = 16'b0000000101000110;
            15'd2133: log10_cal = 16'b0000000101000110;
            15'd2134: log10_cal = 16'b0000000101000110;
            15'd2135: log10_cal = 16'b0000000101000110;
            15'd2136: log10_cal = 16'b0000000101000110;
            15'd2137: log10_cal = 16'b0000000101000111;
            15'd2138: log10_cal = 16'b0000000101000111;
            15'd2139: log10_cal = 16'b0000000101000111;
            15'd2140: log10_cal = 16'b0000000101000111;
            15'd2141: log10_cal = 16'b0000000101001000;
            15'd2142: log10_cal = 16'b0000000101001000;
            15'd2143: log10_cal = 16'b0000000101001000;
            15'd2144: log10_cal = 16'b0000000101001000;
            15'd2145: log10_cal = 16'b0000000101001000;
            15'd2146: log10_cal = 16'b0000000101001001;
            15'd2147: log10_cal = 16'b0000000101001001;
            15'd2148: log10_cal = 16'b0000000101001001;
            15'd2149: log10_cal = 16'b0000000101001001;
            15'd2150: log10_cal = 16'b0000000101001001;
            15'd2151: log10_cal = 16'b0000000101001010;
            15'd2152: log10_cal = 16'b0000000101001010;
            15'd2153: log10_cal = 16'b0000000101001010;
            15'd2154: log10_cal = 16'b0000000101001010;
            15'd2155: log10_cal = 16'b0000000101001010;
            15'd2156: log10_cal = 16'b0000000101001011;
            15'd2157: log10_cal = 16'b0000000101001011;
            15'd2158: log10_cal = 16'b0000000101001011;
            15'd2159: log10_cal = 16'b0000000101001011;
            15'd2160: log10_cal = 16'b0000000101001011;
            15'd2161: log10_cal = 16'b0000000101001100;
            15'd2162: log10_cal = 16'b0000000101001100;
            15'd2163: log10_cal = 16'b0000000101001100;
            15'd2164: log10_cal = 16'b0000000101001100;
            15'd2165: log10_cal = 16'b0000000101001100;
            15'd2166: log10_cal = 16'b0000000101001101;
            15'd2167: log10_cal = 16'b0000000101001101;
            15'd2168: log10_cal = 16'b0000000101001101;
            15'd2169: log10_cal = 16'b0000000101001101;
            15'd2170: log10_cal = 16'b0000000101001101;
            15'd2171: log10_cal = 16'b0000000101001110;
            15'd2172: log10_cal = 16'b0000000101001110;
            15'd2173: log10_cal = 16'b0000000101001110;
            15'd2174: log10_cal = 16'b0000000101001110;
            15'd2175: log10_cal = 16'b0000000101001111;
            15'd2176: log10_cal = 16'b0000000101001111;
            15'd2177: log10_cal = 16'b0000000101001111;
            15'd2178: log10_cal = 16'b0000000101001111;
            15'd2179: log10_cal = 16'b0000000101001111;
            15'd2180: log10_cal = 16'b0000000101010000;
            15'd2181: log10_cal = 16'b0000000101010000;
            15'd2182: log10_cal = 16'b0000000101010000;
            15'd2183: log10_cal = 16'b0000000101010000;
            15'd2184: log10_cal = 16'b0000000101010000;
            15'd2185: log10_cal = 16'b0000000101010001;
            15'd2186: log10_cal = 16'b0000000101010001;
            15'd2187: log10_cal = 16'b0000000101010001;
            15'd2188: log10_cal = 16'b0000000101010001;
            15'd2189: log10_cal = 16'b0000000101010001;
            15'd2190: log10_cal = 16'b0000000101010010;
            15'd2191: log10_cal = 16'b0000000101010010;
            15'd2192: log10_cal = 16'b0000000101010010;
            15'd2193: log10_cal = 16'b0000000101010010;
            15'd2194: log10_cal = 16'b0000000101010010;
            15'd2195: log10_cal = 16'b0000000101010011;
            15'd2196: log10_cal = 16'b0000000101010011;
            15'd2197: log10_cal = 16'b0000000101010011;
            15'd2198: log10_cal = 16'b0000000101010011;
            15'd2199: log10_cal = 16'b0000000101010011;
            15'd2200: log10_cal = 16'b0000000101010100;
            15'd2201: log10_cal = 16'b0000000101010100;
            15'd2202: log10_cal = 16'b0000000101010100;
            15'd2203: log10_cal = 16'b0000000101010100;
            15'd2204: log10_cal = 16'b0000000101010100;
            15'd2205: log10_cal = 16'b0000000101010101;
            15'd2206: log10_cal = 16'b0000000101010101;
            15'd2207: log10_cal = 16'b0000000101010101;
            15'd2208: log10_cal = 16'b0000000101010101;
            15'd2209: log10_cal = 16'b0000000101010101;
            15'd2210: log10_cal = 16'b0000000101010110;
            15'd2211: log10_cal = 16'b0000000101010110;
            15'd2212: log10_cal = 16'b0000000101010110;
            15'd2213: log10_cal = 16'b0000000101010110;
            15'd2214: log10_cal = 16'b0000000101010110;
            15'd2215: log10_cal = 16'b0000000101010111;
            15'd2216: log10_cal = 16'b0000000101010111;
            15'd2217: log10_cal = 16'b0000000101010111;
            15'd2218: log10_cal = 16'b0000000101010111;
            15'd2219: log10_cal = 16'b0000000101010111;
            15'd2220: log10_cal = 16'b0000000101011000;
            15'd2221: log10_cal = 16'b0000000101011000;
            15'd2222: log10_cal = 16'b0000000101011000;
            15'd2223: log10_cal = 16'b0000000101011000;
            15'd2224: log10_cal = 16'b0000000101011000;
            15'd2225: log10_cal = 16'b0000000101011001;
            15'd2226: log10_cal = 16'b0000000101011001;
            15'd2227: log10_cal = 16'b0000000101011001;
            15'd2228: log10_cal = 16'b0000000101011001;
            15'd2229: log10_cal = 16'b0000000101011001;
            15'd2230: log10_cal = 16'b0000000101011010;
            15'd2231: log10_cal = 16'b0000000101011010;
            15'd2232: log10_cal = 16'b0000000101011010;
            15'd2233: log10_cal = 16'b0000000101011010;
            15'd2234: log10_cal = 16'b0000000101011010;
            15'd2235: log10_cal = 16'b0000000101011011;
            15'd2236: log10_cal = 16'b0000000101011011;
            15'd2237: log10_cal = 16'b0000000101011011;
            15'd2238: log10_cal = 16'b0000000101011011;
            15'd2239: log10_cal = 16'b0000000101011011;
            15'd2240: log10_cal = 16'b0000000101011100;
            15'd2241: log10_cal = 16'b0000000101011100;
            15'd2242: log10_cal = 16'b0000000101011100;
            15'd2243: log10_cal = 16'b0000000101011100;
            15'd2244: log10_cal = 16'b0000000101011100;
            15'd2245: log10_cal = 16'b0000000101011101;
            15'd2246: log10_cal = 16'b0000000101011101;
            15'd2247: log10_cal = 16'b0000000101011101;
            15'd2248: log10_cal = 16'b0000000101011101;
            15'd2249: log10_cal = 16'b0000000101011101;
            15'd2250: log10_cal = 16'b0000000101011110;
            15'd2251: log10_cal = 16'b0000000101011110;
            15'd2252: log10_cal = 16'b0000000101011110;
            15'd2253: log10_cal = 16'b0000000101011110;
            15'd2254: log10_cal = 16'b0000000101011110;
            15'd2255: log10_cal = 16'b0000000101011111;
            15'd2256: log10_cal = 16'b0000000101011111;
            15'd2257: log10_cal = 16'b0000000101011111;
            15'd2258: log10_cal = 16'b0000000101011111;
            15'd2259: log10_cal = 16'b0000000101011111;
            15'd2260: log10_cal = 16'b0000000101100000;
            15'd2261: log10_cal = 16'b0000000101100000;
            15'd2262: log10_cal = 16'b0000000101100000;
            15'd2263: log10_cal = 16'b0000000101100000;
            15'd2264: log10_cal = 16'b0000000101100000;
            15'd2265: log10_cal = 16'b0000000101100001;
            15'd2266: log10_cal = 16'b0000000101100001;
            15'd2267: log10_cal = 16'b0000000101100001;
            15'd2268: log10_cal = 16'b0000000101100001;
            15'd2269: log10_cal = 16'b0000000101100001;
            15'd2270: log10_cal = 16'b0000000101100010;
            15'd2271: log10_cal = 16'b0000000101100010;
            15'd2272: log10_cal = 16'b0000000101100010;
            15'd2273: log10_cal = 16'b0000000101100010;
            15'd2274: log10_cal = 16'b0000000101100010;
            15'd2275: log10_cal = 16'b0000000101100011;
            15'd2276: log10_cal = 16'b0000000101100011;
            15'd2277: log10_cal = 16'b0000000101100011;
            15'd2278: log10_cal = 16'b0000000101100011;
            15'd2279: log10_cal = 16'b0000000101100011;
            15'd2280: log10_cal = 16'b0000000101100011;
            15'd2281: log10_cal = 16'b0000000101100100;
            15'd2282: log10_cal = 16'b0000000101100100;
            15'd2283: log10_cal = 16'b0000000101100100;
            15'd2284: log10_cal = 16'b0000000101100100;
            15'd2285: log10_cal = 16'b0000000101100100;
            15'd2286: log10_cal = 16'b0000000101100101;
            15'd2287: log10_cal = 16'b0000000101100101;
            15'd2288: log10_cal = 16'b0000000101100101;
            15'd2289: log10_cal = 16'b0000000101100101;
            15'd2290: log10_cal = 16'b0000000101100101;
            15'd2291: log10_cal = 16'b0000000101100110;
            15'd2292: log10_cal = 16'b0000000101100110;
            15'd2293: log10_cal = 16'b0000000101100110;
            15'd2294: log10_cal = 16'b0000000101100110;
            15'd2295: log10_cal = 16'b0000000101100110;
            15'd2296: log10_cal = 16'b0000000101100111;
            15'd2297: log10_cal = 16'b0000000101100111;
            15'd2298: log10_cal = 16'b0000000101100111;
            15'd2299: log10_cal = 16'b0000000101100111;
            15'd2300: log10_cal = 16'b0000000101100111;
            15'd2301: log10_cal = 16'b0000000101101000;
            15'd2302: log10_cal = 16'b0000000101101000;
            15'd2303: log10_cal = 16'b0000000101101000;
            15'd2304: log10_cal = 16'b0000000101101000;
            15'd2305: log10_cal = 16'b0000000101101000;
            15'd2306: log10_cal = 16'b0000000101101001;
            15'd2307: log10_cal = 16'b0000000101101001;
            15'd2308: log10_cal = 16'b0000000101101001;
            15'd2309: log10_cal = 16'b0000000101101001;
            15'd2310: log10_cal = 16'b0000000101101001;
            15'd2311: log10_cal = 16'b0000000101101001;
            15'd2312: log10_cal = 16'b0000000101101010;
            15'd2313: log10_cal = 16'b0000000101101010;
            15'd2314: log10_cal = 16'b0000000101101010;
            15'd2315: log10_cal = 16'b0000000101101010;
            15'd2316: log10_cal = 16'b0000000101101010;
            15'd2317: log10_cal = 16'b0000000101101011;
            15'd2318: log10_cal = 16'b0000000101101011;
            15'd2319: log10_cal = 16'b0000000101101011;
            15'd2320: log10_cal = 16'b0000000101101011;
            15'd2321: log10_cal = 16'b0000000101101011;
            15'd2322: log10_cal = 16'b0000000101101100;
            15'd2323: log10_cal = 16'b0000000101101100;
            15'd2324: log10_cal = 16'b0000000101101100;
            15'd2325: log10_cal = 16'b0000000101101100;
            15'd2326: log10_cal = 16'b0000000101101100;
            15'd2327: log10_cal = 16'b0000000101101101;
            15'd2328: log10_cal = 16'b0000000101101101;
            15'd2329: log10_cal = 16'b0000000101101101;
            15'd2330: log10_cal = 16'b0000000101101101;
            15'd2331: log10_cal = 16'b0000000101101101;
            15'd2332: log10_cal = 16'b0000000101101110;
            15'd2333: log10_cal = 16'b0000000101101110;
            15'd2334: log10_cal = 16'b0000000101101110;
            15'd2335: log10_cal = 16'b0000000101101110;
            15'd2336: log10_cal = 16'b0000000101101110;
            15'd2337: log10_cal = 16'b0000000101101110;
            15'd2338: log10_cal = 16'b0000000101101111;
            15'd2339: log10_cal = 16'b0000000101101111;
            15'd2340: log10_cal = 16'b0000000101101111;
            15'd2341: log10_cal = 16'b0000000101101111;
            15'd2342: log10_cal = 16'b0000000101101111;
            15'd2343: log10_cal = 16'b0000000101110000;
            15'd2344: log10_cal = 16'b0000000101110000;
            15'd2345: log10_cal = 16'b0000000101110000;
            15'd2346: log10_cal = 16'b0000000101110000;
            15'd2347: log10_cal = 16'b0000000101110000;
            15'd2348: log10_cal = 16'b0000000101110001;
            15'd2349: log10_cal = 16'b0000000101110001;
            15'd2350: log10_cal = 16'b0000000101110001;
            15'd2351: log10_cal = 16'b0000000101110001;
            15'd2352: log10_cal = 16'b0000000101110001;
            15'd2353: log10_cal = 16'b0000000101110001;
            15'd2354: log10_cal = 16'b0000000101110010;
            15'd2355: log10_cal = 16'b0000000101110010;
            15'd2356: log10_cal = 16'b0000000101110010;
            15'd2357: log10_cal = 16'b0000000101110010;
            15'd2358: log10_cal = 16'b0000000101110010;
            15'd2359: log10_cal = 16'b0000000101110011;
            15'd2360: log10_cal = 16'b0000000101110011;
            15'd2361: log10_cal = 16'b0000000101110011;
            15'd2362: log10_cal = 16'b0000000101110011;
            15'd2363: log10_cal = 16'b0000000101110011;
            15'd2364: log10_cal = 16'b0000000101110100;
            15'd2365: log10_cal = 16'b0000000101110100;
            15'd2366: log10_cal = 16'b0000000101110100;
            15'd2367: log10_cal = 16'b0000000101110100;
            15'd2368: log10_cal = 16'b0000000101110100;
            15'd2369: log10_cal = 16'b0000000101110101;
            15'd2370: log10_cal = 16'b0000000101110101;
            15'd2371: log10_cal = 16'b0000000101110101;
            15'd2372: log10_cal = 16'b0000000101110101;
            15'd2373: log10_cal = 16'b0000000101110101;
            15'd2374: log10_cal = 16'b0000000101110101;
            15'd2375: log10_cal = 16'b0000000101110110;
            15'd2376: log10_cal = 16'b0000000101110110;
            15'd2377: log10_cal = 16'b0000000101110110;
            15'd2378: log10_cal = 16'b0000000101110110;
            15'd2379: log10_cal = 16'b0000000101110110;
            15'd2380: log10_cal = 16'b0000000101110111;
            15'd2381: log10_cal = 16'b0000000101110111;
            15'd2382: log10_cal = 16'b0000000101110111;
            15'd2383: log10_cal = 16'b0000000101110111;
            15'd2384: log10_cal = 16'b0000000101110111;
            15'd2385: log10_cal = 16'b0000000101111000;
            15'd2386: log10_cal = 16'b0000000101111000;
            15'd2387: log10_cal = 16'b0000000101111000;
            15'd2388: log10_cal = 16'b0000000101111000;
            15'd2389: log10_cal = 16'b0000000101111000;
            15'd2390: log10_cal = 16'b0000000101111000;
            15'd2391: log10_cal = 16'b0000000101111001;
            15'd2392: log10_cal = 16'b0000000101111001;
            15'd2393: log10_cal = 16'b0000000101111001;
            15'd2394: log10_cal = 16'b0000000101111001;
            15'd2395: log10_cal = 16'b0000000101111001;
            15'd2396: log10_cal = 16'b0000000101111010;
            15'd2397: log10_cal = 16'b0000000101111010;
            15'd2398: log10_cal = 16'b0000000101111010;
            15'd2399: log10_cal = 16'b0000000101111010;
            15'd2400: log10_cal = 16'b0000000101111010;
            15'd2401: log10_cal = 16'b0000000101111010;
            15'd2402: log10_cal = 16'b0000000101111011;
            15'd2403: log10_cal = 16'b0000000101111011;
            15'd2404: log10_cal = 16'b0000000101111011;
            15'd2405: log10_cal = 16'b0000000101111011;
            15'd2406: log10_cal = 16'b0000000101111011;
            15'd2407: log10_cal = 16'b0000000101111100;
            15'd2408: log10_cal = 16'b0000000101111100;
            15'd2409: log10_cal = 16'b0000000101111100;
            15'd2410: log10_cal = 16'b0000000101111100;
            15'd2411: log10_cal = 16'b0000000101111100;
            15'd2412: log10_cal = 16'b0000000101111101;
            15'd2413: log10_cal = 16'b0000000101111101;
            15'd2414: log10_cal = 16'b0000000101111101;
            15'd2415: log10_cal = 16'b0000000101111101;
            15'd2416: log10_cal = 16'b0000000101111101;
            15'd2417: log10_cal = 16'b0000000101111101;
            15'd2418: log10_cal = 16'b0000000101111110;
            15'd2419: log10_cal = 16'b0000000101111110;
            15'd2420: log10_cal = 16'b0000000101111110;
            15'd2421: log10_cal = 16'b0000000101111110;
            15'd2422: log10_cal = 16'b0000000101111110;
            15'd2423: log10_cal = 16'b0000000101111111;
            15'd2424: log10_cal = 16'b0000000101111111;
            15'd2425: log10_cal = 16'b0000000101111111;
            15'd2426: log10_cal = 16'b0000000101111111;
            15'd2427: log10_cal = 16'b0000000101111111;
            15'd2428: log10_cal = 16'b0000000101111111;
            15'd2429: log10_cal = 16'b0000000110000000;
            15'd2430: log10_cal = 16'b0000000110000000;
            15'd2431: log10_cal = 16'b0000000110000000;
            15'd2432: log10_cal = 16'b0000000110000000;
            15'd2433: log10_cal = 16'b0000000110000000;
            15'd2434: log10_cal = 16'b0000000110000001;
            15'd2435: log10_cal = 16'b0000000110000001;
            15'd2436: log10_cal = 16'b0000000110000001;
            15'd2437: log10_cal = 16'b0000000110000001;
            15'd2438: log10_cal = 16'b0000000110000001;
            15'd2439: log10_cal = 16'b0000000110000001;
            15'd2440: log10_cal = 16'b0000000110000010;
            15'd2441: log10_cal = 16'b0000000110000010;
            15'd2442: log10_cal = 16'b0000000110000010;
            15'd2443: log10_cal = 16'b0000000110000010;
            15'd2444: log10_cal = 16'b0000000110000010;
            15'd2445: log10_cal = 16'b0000000110000011;
            15'd2446: log10_cal = 16'b0000000110000011;
            15'd2447: log10_cal = 16'b0000000110000011;
            15'd2448: log10_cal = 16'b0000000110000011;
            15'd2449: log10_cal = 16'b0000000110000011;
            15'd2450: log10_cal = 16'b0000000110000011;
            15'd2451: log10_cal = 16'b0000000110000100;
            15'd2452: log10_cal = 16'b0000000110000100;
            15'd2453: log10_cal = 16'b0000000110000100;
            15'd2454: log10_cal = 16'b0000000110000100;
            15'd2455: log10_cal = 16'b0000000110000100;
            15'd2456: log10_cal = 16'b0000000110000101;
            15'd2457: log10_cal = 16'b0000000110000101;
            15'd2458: log10_cal = 16'b0000000110000101;
            15'd2459: log10_cal = 16'b0000000110000101;
            15'd2460: log10_cal = 16'b0000000110000101;
            15'd2461: log10_cal = 16'b0000000110000101;
            15'd2462: log10_cal = 16'b0000000110000110;
            15'd2463: log10_cal = 16'b0000000110000110;
            15'd2464: log10_cal = 16'b0000000110000110;
            15'd2465: log10_cal = 16'b0000000110000110;
            15'd2466: log10_cal = 16'b0000000110000110;
            15'd2467: log10_cal = 16'b0000000110000111;
            15'd2468: log10_cal = 16'b0000000110000111;
            15'd2469: log10_cal = 16'b0000000110000111;
            15'd2470: log10_cal = 16'b0000000110000111;
            15'd2471: log10_cal = 16'b0000000110000111;
            15'd2472: log10_cal = 16'b0000000110000111;
            15'd2473: log10_cal = 16'b0000000110001000;
            15'd2474: log10_cal = 16'b0000000110001000;
            15'd2475: log10_cal = 16'b0000000110001000;
            15'd2476: log10_cal = 16'b0000000110001000;
            15'd2477: log10_cal = 16'b0000000110001000;
            15'd2478: log10_cal = 16'b0000000110001001;
            15'd2479: log10_cal = 16'b0000000110001001;
            15'd2480: log10_cal = 16'b0000000110001001;
            15'd2481: log10_cal = 16'b0000000110001001;
            15'd2482: log10_cal = 16'b0000000110001001;
            15'd2483: log10_cal = 16'b0000000110001001;
            15'd2484: log10_cal = 16'b0000000110001010;
            15'd2485: log10_cal = 16'b0000000110001010;
            15'd2486: log10_cal = 16'b0000000110001010;
            15'd2487: log10_cal = 16'b0000000110001010;
            15'd2488: log10_cal = 16'b0000000110001010;
            15'd2489: log10_cal = 16'b0000000110001010;
            15'd2490: log10_cal = 16'b0000000110001011;
            15'd2491: log10_cal = 16'b0000000110001011;
            15'd2492: log10_cal = 16'b0000000110001011;
            15'd2493: log10_cal = 16'b0000000110001011;
            15'd2494: log10_cal = 16'b0000000110001011;
            15'd2495: log10_cal = 16'b0000000110001100;
            15'd2496: log10_cal = 16'b0000000110001100;
            15'd2497: log10_cal = 16'b0000000110001100;
            15'd2498: log10_cal = 16'b0000000110001100;
            15'd2499: log10_cal = 16'b0000000110001100;
            15'd2500: log10_cal = 16'b0000000110001100;
            15'd2501: log10_cal = 16'b0000000110001101;
            15'd2502: log10_cal = 16'b0000000110001101;
            15'd2503: log10_cal = 16'b0000000110001101;
            15'd2504: log10_cal = 16'b0000000110001101;
            15'd2505: log10_cal = 16'b0000000110001101;
            15'd2506: log10_cal = 16'b0000000110001110;
            15'd2507: log10_cal = 16'b0000000110001110;
            15'd2508: log10_cal = 16'b0000000110001110;
            15'd2509: log10_cal = 16'b0000000110001110;
            15'd2510: log10_cal = 16'b0000000110001110;
            15'd2511: log10_cal = 16'b0000000110001110;
            15'd2512: log10_cal = 16'b0000000110001111;
            15'd2513: log10_cal = 16'b0000000110001111;
            15'd2514: log10_cal = 16'b0000000110001111;
            15'd2515: log10_cal = 16'b0000000110001111;
            15'd2516: log10_cal = 16'b0000000110001111;
            15'd2517: log10_cal = 16'b0000000110001111;
            15'd2518: log10_cal = 16'b0000000110010000;
            15'd2519: log10_cal = 16'b0000000110010000;
            15'd2520: log10_cal = 16'b0000000110010000;
            15'd2521: log10_cal = 16'b0000000110010000;
            15'd2522: log10_cal = 16'b0000000110010000;
            15'd2523: log10_cal = 16'b0000000110010001;
            15'd2524: log10_cal = 16'b0000000110010001;
            15'd2525: log10_cal = 16'b0000000110010001;
            15'd2526: log10_cal = 16'b0000000110010001;
            15'd2527: log10_cal = 16'b0000000110010001;
            15'd2528: log10_cal = 16'b0000000110010001;
            15'd2529: log10_cal = 16'b0000000110010010;
            15'd2530: log10_cal = 16'b0000000110010010;
            15'd2531: log10_cal = 16'b0000000110010010;
            15'd2532: log10_cal = 16'b0000000110010010;
            15'd2533: log10_cal = 16'b0000000110010010;
            15'd2534: log10_cal = 16'b0000000110010010;
            15'd2535: log10_cal = 16'b0000000110010011;
            15'd2536: log10_cal = 16'b0000000110010011;
            15'd2537: log10_cal = 16'b0000000110010011;
            15'd2538: log10_cal = 16'b0000000110010011;
            15'd2539: log10_cal = 16'b0000000110010011;
            15'd2540: log10_cal = 16'b0000000110010100;
            15'd2541: log10_cal = 16'b0000000110010100;
            15'd2542: log10_cal = 16'b0000000110010100;
            15'd2543: log10_cal = 16'b0000000110010100;
            15'd2544: log10_cal = 16'b0000000110010100;
            15'd2545: log10_cal = 16'b0000000110010100;
            15'd2546: log10_cal = 16'b0000000110010101;
            15'd2547: log10_cal = 16'b0000000110010101;
            15'd2548: log10_cal = 16'b0000000110010101;
            15'd2549: log10_cal = 16'b0000000110010101;
            15'd2550: log10_cal = 16'b0000000110010101;
            15'd2551: log10_cal = 16'b0000000110010101;
            15'd2552: log10_cal = 16'b0000000110010110;
            15'd2553: log10_cal = 16'b0000000110010110;
            15'd2554: log10_cal = 16'b0000000110010110;
            15'd2555: log10_cal = 16'b0000000110010110;
            15'd2556: log10_cal = 16'b0000000110010110;
            15'd2557: log10_cal = 16'b0000000110010110;
            15'd2558: log10_cal = 16'b0000000110010111;
            15'd2559: log10_cal = 16'b0000000110010111;
            15'd2560: log10_cal = 16'b0000000110010111;
            15'd2561: log10_cal = 16'b0000000110010111;
            15'd2562: log10_cal = 16'b0000000110010111;
            15'd2563: log10_cal = 16'b0000000110011000;
            15'd2564: log10_cal = 16'b0000000110011000;
            15'd2565: log10_cal = 16'b0000000110011000;
            15'd2566: log10_cal = 16'b0000000110011000;
            15'd2567: log10_cal = 16'b0000000110011000;
            15'd2568: log10_cal = 16'b0000000110011000;
            15'd2569: log10_cal = 16'b0000000110011001;
            15'd2570: log10_cal = 16'b0000000110011001;
            15'd2571: log10_cal = 16'b0000000110011001;
            15'd2572: log10_cal = 16'b0000000110011001;
            15'd2573: log10_cal = 16'b0000000110011001;
            15'd2574: log10_cal = 16'b0000000110011001;
            15'd2575: log10_cal = 16'b0000000110011010;
            15'd2576: log10_cal = 16'b0000000110011010;
            15'd2577: log10_cal = 16'b0000000110011010;
            15'd2578: log10_cal = 16'b0000000110011010;
            15'd2579: log10_cal = 16'b0000000110011010;
            15'd2580: log10_cal = 16'b0000000110011010;
            15'd2581: log10_cal = 16'b0000000110011011;
            15'd2582: log10_cal = 16'b0000000110011011;
            15'd2583: log10_cal = 16'b0000000110011011;
            15'd2584: log10_cal = 16'b0000000110011011;
            15'd2585: log10_cal = 16'b0000000110011011;
            15'd2586: log10_cal = 16'b0000000110011011;
            15'd2587: log10_cal = 16'b0000000110011100;
            15'd2588: log10_cal = 16'b0000000110011100;
            15'd2589: log10_cal = 16'b0000000110011100;
            15'd2590: log10_cal = 16'b0000000110011100;
            15'd2591: log10_cal = 16'b0000000110011100;
            15'd2592: log10_cal = 16'b0000000110011101;
            15'd2593: log10_cal = 16'b0000000110011101;
            15'd2594: log10_cal = 16'b0000000110011101;
            15'd2595: log10_cal = 16'b0000000110011101;
            15'd2596: log10_cal = 16'b0000000110011101;
            15'd2597: log10_cal = 16'b0000000110011101;
            15'd2598: log10_cal = 16'b0000000110011110;
            15'd2599: log10_cal = 16'b0000000110011110;
            15'd2600: log10_cal = 16'b0000000110011110;
            15'd2601: log10_cal = 16'b0000000110011110;
            15'd2602: log10_cal = 16'b0000000110011110;
            15'd2603: log10_cal = 16'b0000000110011110;
            15'd2604: log10_cal = 16'b0000000110011111;
            15'd2605: log10_cal = 16'b0000000110011111;
            15'd2606: log10_cal = 16'b0000000110011111;
            15'd2607: log10_cal = 16'b0000000110011111;
            15'd2608: log10_cal = 16'b0000000110011111;
            15'd2609: log10_cal = 16'b0000000110011111;
            15'd2610: log10_cal = 16'b0000000110100000;
            15'd2611: log10_cal = 16'b0000000110100000;
            15'd2612: log10_cal = 16'b0000000110100000;
            15'd2613: log10_cal = 16'b0000000110100000;
            15'd2614: log10_cal = 16'b0000000110100000;
            15'd2615: log10_cal = 16'b0000000110100000;
            15'd2616: log10_cal = 16'b0000000110100001;
            15'd2617: log10_cal = 16'b0000000110100001;
            15'd2618: log10_cal = 16'b0000000110100001;
            15'd2619: log10_cal = 16'b0000000110100001;
            15'd2620: log10_cal = 16'b0000000110100001;
            15'd2621: log10_cal = 16'b0000000110100001;
            15'd2622: log10_cal = 16'b0000000110100010;
            15'd2623: log10_cal = 16'b0000000110100010;
            15'd2624: log10_cal = 16'b0000000110100010;
            15'd2625: log10_cal = 16'b0000000110100010;
            15'd2626: log10_cal = 16'b0000000110100010;
            15'd2627: log10_cal = 16'b0000000110100010;
            15'd2628: log10_cal = 16'b0000000110100011;
            15'd2629: log10_cal = 16'b0000000110100011;
            15'd2630: log10_cal = 16'b0000000110100011;
            15'd2631: log10_cal = 16'b0000000110100011;
            15'd2632: log10_cal = 16'b0000000110100011;
            15'd2633: log10_cal = 16'b0000000110100011;
            15'd2634: log10_cal = 16'b0000000110100100;
            15'd2635: log10_cal = 16'b0000000110100100;
            15'd2636: log10_cal = 16'b0000000110100100;
            15'd2637: log10_cal = 16'b0000000110100100;
            15'd2638: log10_cal = 16'b0000000110100100;
            15'd2639: log10_cal = 16'b0000000110100101;
            15'd2640: log10_cal = 16'b0000000110100101;
            15'd2641: log10_cal = 16'b0000000110100101;
            15'd2642: log10_cal = 16'b0000000110100101;
            15'd2643: log10_cal = 16'b0000000110100101;
            15'd2644: log10_cal = 16'b0000000110100101;
            15'd2645: log10_cal = 16'b0000000110100110;
            15'd2646: log10_cal = 16'b0000000110100110;
            15'd2647: log10_cal = 16'b0000000110100110;
            15'd2648: log10_cal = 16'b0000000110100110;
            15'd2649: log10_cal = 16'b0000000110100110;
            15'd2650: log10_cal = 16'b0000000110100110;
            15'd2651: log10_cal = 16'b0000000110100111;
            15'd2652: log10_cal = 16'b0000000110100111;
            15'd2653: log10_cal = 16'b0000000110100111;
            15'd2654: log10_cal = 16'b0000000110100111;
            15'd2655: log10_cal = 16'b0000000110100111;
            15'd2656: log10_cal = 16'b0000000110100111;
            15'd2657: log10_cal = 16'b0000000110101000;
            15'd2658: log10_cal = 16'b0000000110101000;
            15'd2659: log10_cal = 16'b0000000110101000;
            15'd2660: log10_cal = 16'b0000000110101000;
            15'd2661: log10_cal = 16'b0000000110101000;
            15'd2662: log10_cal = 16'b0000000110101000;
            15'd2663: log10_cal = 16'b0000000110101001;
            15'd2664: log10_cal = 16'b0000000110101001;
            15'd2665: log10_cal = 16'b0000000110101001;
            15'd2666: log10_cal = 16'b0000000110101001;
            15'd2667: log10_cal = 16'b0000000110101001;
            15'd2668: log10_cal = 16'b0000000110101001;
            15'd2669: log10_cal = 16'b0000000110101010;
            15'd2670: log10_cal = 16'b0000000110101010;
            15'd2671: log10_cal = 16'b0000000110101010;
            15'd2672: log10_cal = 16'b0000000110101010;
            15'd2673: log10_cal = 16'b0000000110101010;
            15'd2674: log10_cal = 16'b0000000110101010;
            15'd2675: log10_cal = 16'b0000000110101011;
            15'd2676: log10_cal = 16'b0000000110101011;
            15'd2677: log10_cal = 16'b0000000110101011;
            15'd2678: log10_cal = 16'b0000000110101011;
            15'd2679: log10_cal = 16'b0000000110101011;
            15'd2680: log10_cal = 16'b0000000110101011;
            15'd2681: log10_cal = 16'b0000000110101100;
            15'd2682: log10_cal = 16'b0000000110101100;
            15'd2683: log10_cal = 16'b0000000110101100;
            15'd2684: log10_cal = 16'b0000000110101100;
            15'd2685: log10_cal = 16'b0000000110101100;
            15'd2686: log10_cal = 16'b0000000110101100;
            15'd2687: log10_cal = 16'b0000000110101101;
            15'd2688: log10_cal = 16'b0000000110101101;
            15'd2689: log10_cal = 16'b0000000110101101;
            15'd2690: log10_cal = 16'b0000000110101101;
            15'd2691: log10_cal = 16'b0000000110101101;
            15'd2692: log10_cal = 16'b0000000110101101;
            15'd2693: log10_cal = 16'b0000000110101110;
            15'd2694: log10_cal = 16'b0000000110101110;
            15'd2695: log10_cal = 16'b0000000110101110;
            15'd2696: log10_cal = 16'b0000000110101110;
            15'd2697: log10_cal = 16'b0000000110101110;
            15'd2698: log10_cal = 16'b0000000110101110;
            15'd2699: log10_cal = 16'b0000000110101111;
            15'd2700: log10_cal = 16'b0000000110101111;
            15'd2701: log10_cal = 16'b0000000110101111;
            15'd2702: log10_cal = 16'b0000000110101111;
            15'd2703: log10_cal = 16'b0000000110101111;
            15'd2704: log10_cal = 16'b0000000110101111;
            15'd2705: log10_cal = 16'b0000000110101111;
            15'd2706: log10_cal = 16'b0000000110110000;
            15'd2707: log10_cal = 16'b0000000110110000;
            15'd2708: log10_cal = 16'b0000000110110000;
            15'd2709: log10_cal = 16'b0000000110110000;
            15'd2710: log10_cal = 16'b0000000110110000;
            15'd2711: log10_cal = 16'b0000000110110000;
            15'd2712: log10_cal = 16'b0000000110110001;
            15'd2713: log10_cal = 16'b0000000110110001;
            15'd2714: log10_cal = 16'b0000000110110001;
            15'd2715: log10_cal = 16'b0000000110110001;
            15'd2716: log10_cal = 16'b0000000110110001;
            15'd2717: log10_cal = 16'b0000000110110001;
            15'd2718: log10_cal = 16'b0000000110110010;
            15'd2719: log10_cal = 16'b0000000110110010;
            15'd2720: log10_cal = 16'b0000000110110010;
            15'd2721: log10_cal = 16'b0000000110110010;
            15'd2722: log10_cal = 16'b0000000110110010;
            15'd2723: log10_cal = 16'b0000000110110010;
            15'd2724: log10_cal = 16'b0000000110110011;
            15'd2725: log10_cal = 16'b0000000110110011;
            15'd2726: log10_cal = 16'b0000000110110011;
            15'd2727: log10_cal = 16'b0000000110110011;
            15'd2728: log10_cal = 16'b0000000110110011;
            15'd2729: log10_cal = 16'b0000000110110011;
            15'd2730: log10_cal = 16'b0000000110110100;
            15'd2731: log10_cal = 16'b0000000110110100;
            15'd2732: log10_cal = 16'b0000000110110100;
            15'd2733: log10_cal = 16'b0000000110110100;
            15'd2734: log10_cal = 16'b0000000110110100;
            15'd2735: log10_cal = 16'b0000000110110100;
            15'd2736: log10_cal = 16'b0000000110110101;
            15'd2737: log10_cal = 16'b0000000110110101;
            15'd2738: log10_cal = 16'b0000000110110101;
            15'd2739: log10_cal = 16'b0000000110110101;
            15'd2740: log10_cal = 16'b0000000110110101;
            15'd2741: log10_cal = 16'b0000000110110101;
            15'd2742: log10_cal = 16'b0000000110110110;
            15'd2743: log10_cal = 16'b0000000110110110;
            15'd2744: log10_cal = 16'b0000000110110110;
            15'd2745: log10_cal = 16'b0000000110110110;
            15'd2746: log10_cal = 16'b0000000110110110;
            15'd2747: log10_cal = 16'b0000000110110110;
            15'd2748: log10_cal = 16'b0000000110110111;
            15'd2749: log10_cal = 16'b0000000110110111;
            15'd2750: log10_cal = 16'b0000000110110111;
            15'd2751: log10_cal = 16'b0000000110110111;
            15'd2752: log10_cal = 16'b0000000110110111;
            15'd2753: log10_cal = 16'b0000000110110111;
            15'd2754: log10_cal = 16'b0000000110110111;
            15'd2755: log10_cal = 16'b0000000110111000;
            15'd2756: log10_cal = 16'b0000000110111000;
            15'd2757: log10_cal = 16'b0000000110111000;
            15'd2758: log10_cal = 16'b0000000110111000;
            15'd2759: log10_cal = 16'b0000000110111000;
            15'd2760: log10_cal = 16'b0000000110111000;
            15'd2761: log10_cal = 16'b0000000110111001;
            15'd2762: log10_cal = 16'b0000000110111001;
            15'd2763: log10_cal = 16'b0000000110111001;
            15'd2764: log10_cal = 16'b0000000110111001;
            15'd2765: log10_cal = 16'b0000000110111001;
            15'd2766: log10_cal = 16'b0000000110111001;
            15'd2767: log10_cal = 16'b0000000110111010;
            15'd2768: log10_cal = 16'b0000000110111010;
            15'd2769: log10_cal = 16'b0000000110111010;
            15'd2770: log10_cal = 16'b0000000110111010;
            15'd2771: log10_cal = 16'b0000000110111010;
            15'd2772: log10_cal = 16'b0000000110111010;
            15'd2773: log10_cal = 16'b0000000110111011;
            15'd2774: log10_cal = 16'b0000000110111011;
            15'd2775: log10_cal = 16'b0000000110111011;
            15'd2776: log10_cal = 16'b0000000110111011;
            15'd2777: log10_cal = 16'b0000000110111011;
            15'd2778: log10_cal = 16'b0000000110111011;
            15'd2779: log10_cal = 16'b0000000110111011;
            15'd2780: log10_cal = 16'b0000000110111100;
            15'd2781: log10_cal = 16'b0000000110111100;
            15'd2782: log10_cal = 16'b0000000110111100;
            15'd2783: log10_cal = 16'b0000000110111100;
            15'd2784: log10_cal = 16'b0000000110111100;
            15'd2785: log10_cal = 16'b0000000110111100;
            15'd2786: log10_cal = 16'b0000000110111101;
            15'd2787: log10_cal = 16'b0000000110111101;
            15'd2788: log10_cal = 16'b0000000110111101;
            15'd2789: log10_cal = 16'b0000000110111101;
            15'd2790: log10_cal = 16'b0000000110111101;
            15'd2791: log10_cal = 16'b0000000110111101;
            15'd2792: log10_cal = 16'b0000000110111110;
            15'd2793: log10_cal = 16'b0000000110111110;
            15'd2794: log10_cal = 16'b0000000110111110;
            15'd2795: log10_cal = 16'b0000000110111110;
            15'd2796: log10_cal = 16'b0000000110111110;
            15'd2797: log10_cal = 16'b0000000110111110;
            15'd2798: log10_cal = 16'b0000000110111111;
            15'd2799: log10_cal = 16'b0000000110111111;
            15'd2800: log10_cal = 16'b0000000110111111;
            15'd2801: log10_cal = 16'b0000000110111111;
            15'd2802: log10_cal = 16'b0000000110111111;
            15'd2803: log10_cal = 16'b0000000110111111;
            15'd2804: log10_cal = 16'b0000000110111111;
            15'd2805: log10_cal = 16'b0000000111000000;
            15'd2806: log10_cal = 16'b0000000111000000;
            15'd2807: log10_cal = 16'b0000000111000000;
            15'd2808: log10_cal = 16'b0000000111000000;
            15'd2809: log10_cal = 16'b0000000111000000;
            15'd2810: log10_cal = 16'b0000000111000000;
            15'd2811: log10_cal = 16'b0000000111000001;
            15'd2812: log10_cal = 16'b0000000111000001;
            15'd2813: log10_cal = 16'b0000000111000001;
            15'd2814: log10_cal = 16'b0000000111000001;
            15'd2815: log10_cal = 16'b0000000111000001;
            15'd2816: log10_cal = 16'b0000000111000001;
            15'd2817: log10_cal = 16'b0000000111000010;
            15'd2818: log10_cal = 16'b0000000111000010;
            15'd2819: log10_cal = 16'b0000000111000010;
            15'd2820: log10_cal = 16'b0000000111000010;
            15'd2821: log10_cal = 16'b0000000111000010;
            15'd2822: log10_cal = 16'b0000000111000010;
            15'd2823: log10_cal = 16'b0000000111000010;
            15'd2824: log10_cal = 16'b0000000111000011;
            15'd2825: log10_cal = 16'b0000000111000011;
            15'd2826: log10_cal = 16'b0000000111000011;
            15'd2827: log10_cal = 16'b0000000111000011;
            15'd2828: log10_cal = 16'b0000000111000011;
            15'd2829: log10_cal = 16'b0000000111000011;
            15'd2830: log10_cal = 16'b0000000111000100;
            15'd2831: log10_cal = 16'b0000000111000100;
            15'd2832: log10_cal = 16'b0000000111000100;
            15'd2833: log10_cal = 16'b0000000111000100;
            15'd2834: log10_cal = 16'b0000000111000100;
            15'd2835: log10_cal = 16'b0000000111000100;
            15'd2836: log10_cal = 16'b0000000111000101;
            15'd2837: log10_cal = 16'b0000000111000101;
            15'd2838: log10_cal = 16'b0000000111000101;
            15'd2839: log10_cal = 16'b0000000111000101;
            15'd2840: log10_cal = 16'b0000000111000101;
            15'd2841: log10_cal = 16'b0000000111000101;
            15'd2842: log10_cal = 16'b0000000111000101;
            15'd2843: log10_cal = 16'b0000000111000110;
            15'd2844: log10_cal = 16'b0000000111000110;
            15'd2845: log10_cal = 16'b0000000111000110;
            15'd2846: log10_cal = 16'b0000000111000110;
            15'd2847: log10_cal = 16'b0000000111000110;
            15'd2848: log10_cal = 16'b0000000111000110;
            15'd2849: log10_cal = 16'b0000000111000111;
            15'd2850: log10_cal = 16'b0000000111000111;
            15'd2851: log10_cal = 16'b0000000111000111;
            15'd2852: log10_cal = 16'b0000000111000111;
            15'd2853: log10_cal = 16'b0000000111000111;
            15'd2854: log10_cal = 16'b0000000111000111;
            15'd2855: log10_cal = 16'b0000000111000111;
            15'd2856: log10_cal = 16'b0000000111001000;
            15'd2857: log10_cal = 16'b0000000111001000;
            15'd2858: log10_cal = 16'b0000000111001000;
            15'd2859: log10_cal = 16'b0000000111001000;
            15'd2860: log10_cal = 16'b0000000111001000;
            15'd2861: log10_cal = 16'b0000000111001000;
            15'd2862: log10_cal = 16'b0000000111001001;
            15'd2863: log10_cal = 16'b0000000111001001;
            15'd2864: log10_cal = 16'b0000000111001001;
            15'd2865: log10_cal = 16'b0000000111001001;
            15'd2866: log10_cal = 16'b0000000111001001;
            15'd2867: log10_cal = 16'b0000000111001001;
            15'd2868: log10_cal = 16'b0000000111001010;
            15'd2869: log10_cal = 16'b0000000111001010;
            15'd2870: log10_cal = 16'b0000000111001010;
            15'd2871: log10_cal = 16'b0000000111001010;
            15'd2872: log10_cal = 16'b0000000111001010;
            15'd2873: log10_cal = 16'b0000000111001010;
            15'd2874: log10_cal = 16'b0000000111001010;
            15'd2875: log10_cal = 16'b0000000111001011;
            15'd2876: log10_cal = 16'b0000000111001011;
            15'd2877: log10_cal = 16'b0000000111001011;
            15'd2878: log10_cal = 16'b0000000111001011;
            15'd2879: log10_cal = 16'b0000000111001011;
            15'd2880: log10_cal = 16'b0000000111001011;
            15'd2881: log10_cal = 16'b0000000111001100;
            15'd2882: log10_cal = 16'b0000000111001100;
            15'd2883: log10_cal = 16'b0000000111001100;
            15'd2884: log10_cal = 16'b0000000111001100;
            15'd2885: log10_cal = 16'b0000000111001100;
            15'd2886: log10_cal = 16'b0000000111001100;
            15'd2887: log10_cal = 16'b0000000111001100;
            15'd2888: log10_cal = 16'b0000000111001101;
            15'd2889: log10_cal = 16'b0000000111001101;
            15'd2890: log10_cal = 16'b0000000111001101;
            15'd2891: log10_cal = 16'b0000000111001101;
            15'd2892: log10_cal = 16'b0000000111001101;
            15'd2893: log10_cal = 16'b0000000111001101;
            15'd2894: log10_cal = 16'b0000000111001110;
            15'd2895: log10_cal = 16'b0000000111001110;
            15'd2896: log10_cal = 16'b0000000111001110;
            15'd2897: log10_cal = 16'b0000000111001110;
            15'd2898: log10_cal = 16'b0000000111001110;
            15'd2899: log10_cal = 16'b0000000111001110;
            15'd2900: log10_cal = 16'b0000000111001110;
            15'd2901: log10_cal = 16'b0000000111001111;
            15'd2902: log10_cal = 16'b0000000111001111;
            15'd2903: log10_cal = 16'b0000000111001111;
            15'd2904: log10_cal = 16'b0000000111001111;
            15'd2905: log10_cal = 16'b0000000111001111;
            15'd2906: log10_cal = 16'b0000000111001111;
            15'd2907: log10_cal = 16'b0000000111010000;
            15'd2908: log10_cal = 16'b0000000111010000;
            15'd2909: log10_cal = 16'b0000000111010000;
            15'd2910: log10_cal = 16'b0000000111010000;
            15'd2911: log10_cal = 16'b0000000111010000;
            15'd2912: log10_cal = 16'b0000000111010000;
            15'd2913: log10_cal = 16'b0000000111010000;
            15'd2914: log10_cal = 16'b0000000111010001;
            15'd2915: log10_cal = 16'b0000000111010001;
            15'd2916: log10_cal = 16'b0000000111010001;
            15'd2917: log10_cal = 16'b0000000111010001;
            15'd2918: log10_cal = 16'b0000000111010001;
            15'd2919: log10_cal = 16'b0000000111010001;
            15'd2920: log10_cal = 16'b0000000111010010;
            15'd2921: log10_cal = 16'b0000000111010010;
            15'd2922: log10_cal = 16'b0000000111010010;
            15'd2923: log10_cal = 16'b0000000111010010;
            15'd2924: log10_cal = 16'b0000000111010010;
            15'd2925: log10_cal = 16'b0000000111010010;
            15'd2926: log10_cal = 16'b0000000111010010;
            15'd2927: log10_cal = 16'b0000000111010011;
            15'd2928: log10_cal = 16'b0000000111010011;
            15'd2929: log10_cal = 16'b0000000111010011;
            15'd2930: log10_cal = 16'b0000000111010011;
            15'd2931: log10_cal = 16'b0000000111010011;
            15'd2932: log10_cal = 16'b0000000111010011;
            15'd2933: log10_cal = 16'b0000000111010011;
            15'd2934: log10_cal = 16'b0000000111010100;
            15'd2935: log10_cal = 16'b0000000111010100;
            15'd2936: log10_cal = 16'b0000000111010100;
            15'd2937: log10_cal = 16'b0000000111010100;
            15'd2938: log10_cal = 16'b0000000111010100;
            15'd2939: log10_cal = 16'b0000000111010100;
            15'd2940: log10_cal = 16'b0000000111010101;
            15'd2941: log10_cal = 16'b0000000111010101;
            15'd2942: log10_cal = 16'b0000000111010101;
            15'd2943: log10_cal = 16'b0000000111010101;
            15'd2944: log10_cal = 16'b0000000111010101;
            15'd2945: log10_cal = 16'b0000000111010101;
            15'd2946: log10_cal = 16'b0000000111010101;
            15'd2947: log10_cal = 16'b0000000111010110;
            15'd2948: log10_cal = 16'b0000000111010110;
            15'd2949: log10_cal = 16'b0000000111010110;
            15'd2950: log10_cal = 16'b0000000111010110;
            15'd2951: log10_cal = 16'b0000000111010110;
            15'd2952: log10_cal = 16'b0000000111010110;
            15'd2953: log10_cal = 16'b0000000111010111;
            15'd2954: log10_cal = 16'b0000000111010111;
            15'd2955: log10_cal = 16'b0000000111010111;
            15'd2956: log10_cal = 16'b0000000111010111;
            15'd2957: log10_cal = 16'b0000000111010111;
            15'd2958: log10_cal = 16'b0000000111010111;
            15'd2959: log10_cal = 16'b0000000111010111;
            15'd2960: log10_cal = 16'b0000000111011000;
            15'd2961: log10_cal = 16'b0000000111011000;
            15'd2962: log10_cal = 16'b0000000111011000;
            15'd2963: log10_cal = 16'b0000000111011000;
            15'd2964: log10_cal = 16'b0000000111011000;
            15'd2965: log10_cal = 16'b0000000111011000;
            15'd2966: log10_cal = 16'b0000000111011000;
            15'd2967: log10_cal = 16'b0000000111011001;
            15'd2968: log10_cal = 16'b0000000111011001;
            15'd2969: log10_cal = 16'b0000000111011001;
            15'd2970: log10_cal = 16'b0000000111011001;
            15'd2971: log10_cal = 16'b0000000111011001;
            15'd2972: log10_cal = 16'b0000000111011001;
            15'd2973: log10_cal = 16'b0000000111011010;
            15'd2974: log10_cal = 16'b0000000111011010;
            15'd2975: log10_cal = 16'b0000000111011010;
            15'd2976: log10_cal = 16'b0000000111011010;
            15'd2977: log10_cal = 16'b0000000111011010;
            15'd2978: log10_cal = 16'b0000000111011010;
            15'd2979: log10_cal = 16'b0000000111011010;
            15'd2980: log10_cal = 16'b0000000111011011;
            15'd2981: log10_cal = 16'b0000000111011011;
            15'd2982: log10_cal = 16'b0000000111011011;
            15'd2983: log10_cal = 16'b0000000111011011;
            15'd2984: log10_cal = 16'b0000000111011011;
            15'd2985: log10_cal = 16'b0000000111011011;
            15'd2986: log10_cal = 16'b0000000111011011;
            15'd2987: log10_cal = 16'b0000000111011100;
            15'd2988: log10_cal = 16'b0000000111011100;
            15'd2989: log10_cal = 16'b0000000111011100;
            15'd2990: log10_cal = 16'b0000000111011100;
            15'd2991: log10_cal = 16'b0000000111011100;
            15'd2992: log10_cal = 16'b0000000111011100;
            15'd2993: log10_cal = 16'b0000000111011100;
            15'd2994: log10_cal = 16'b0000000111011101;
            15'd2995: log10_cal = 16'b0000000111011101;
            15'd2996: log10_cal = 16'b0000000111011101;
            15'd2997: log10_cal = 16'b0000000111011101;
            15'd2998: log10_cal = 16'b0000000111011101;
            15'd2999: log10_cal = 16'b0000000111011101;
            15'd3000: log10_cal = 16'b0000000111011110;
            15'd3001: log10_cal = 16'b0000000111011110;
            15'd3002: log10_cal = 16'b0000000111011110;
            15'd3003: log10_cal = 16'b0000000111011110;
            15'd3004: log10_cal = 16'b0000000111011110;
            15'd3005: log10_cal = 16'b0000000111011110;
            15'd3006: log10_cal = 16'b0000000111011110;
            15'd3007: log10_cal = 16'b0000000111011111;
            15'd3008: log10_cal = 16'b0000000111011111;
            15'd3009: log10_cal = 16'b0000000111011111;
            15'd3010: log10_cal = 16'b0000000111011111;
            15'd3011: log10_cal = 16'b0000000111011111;
            15'd3012: log10_cal = 16'b0000000111011111;
            15'd3013: log10_cal = 16'b0000000111011111;
            15'd3014: log10_cal = 16'b0000000111100000;
            15'd3015: log10_cal = 16'b0000000111100000;
            15'd3016: log10_cal = 16'b0000000111100000;
            15'd3017: log10_cal = 16'b0000000111100000;
            15'd3018: log10_cal = 16'b0000000111100000;
            15'd3019: log10_cal = 16'b0000000111100000;
            15'd3020: log10_cal = 16'b0000000111100000;
            15'd3021: log10_cal = 16'b0000000111100001;
            15'd3022: log10_cal = 16'b0000000111100001;
            15'd3023: log10_cal = 16'b0000000111100001;
            15'd3024: log10_cal = 16'b0000000111100001;
            15'd3025: log10_cal = 16'b0000000111100001;
            15'd3026: log10_cal = 16'b0000000111100001;
            15'd3027: log10_cal = 16'b0000000111100010;
            15'd3028: log10_cal = 16'b0000000111100010;
            15'd3029: log10_cal = 16'b0000000111100010;
            15'd3030: log10_cal = 16'b0000000111100010;
            15'd3031: log10_cal = 16'b0000000111100010;
            15'd3032: log10_cal = 16'b0000000111100010;
            15'd3033: log10_cal = 16'b0000000111100010;
            15'd3034: log10_cal = 16'b0000000111100011;
            15'd3035: log10_cal = 16'b0000000111100011;
            15'd3036: log10_cal = 16'b0000000111100011;
            15'd3037: log10_cal = 16'b0000000111100011;
            15'd3038: log10_cal = 16'b0000000111100011;
            15'd3039: log10_cal = 16'b0000000111100011;
            15'd3040: log10_cal = 16'b0000000111100011;
            15'd3041: log10_cal = 16'b0000000111100100;
            15'd3042: log10_cal = 16'b0000000111100100;
            15'd3043: log10_cal = 16'b0000000111100100;
            15'd3044: log10_cal = 16'b0000000111100100;
            15'd3045: log10_cal = 16'b0000000111100100;
            15'd3046: log10_cal = 16'b0000000111100100;
            15'd3047: log10_cal = 16'b0000000111100100;
            15'd3048: log10_cal = 16'b0000000111100101;
            15'd3049: log10_cal = 16'b0000000111100101;
            15'd3050: log10_cal = 16'b0000000111100101;
            15'd3051: log10_cal = 16'b0000000111100101;
            15'd3052: log10_cal = 16'b0000000111100101;
            15'd3053: log10_cal = 16'b0000000111100101;
            15'd3054: log10_cal = 16'b0000000111100101;
            15'd3055: log10_cal = 16'b0000000111100110;
            15'd3056: log10_cal = 16'b0000000111100110;
            15'd3057: log10_cal = 16'b0000000111100110;
            15'd3058: log10_cal = 16'b0000000111100110;
            15'd3059: log10_cal = 16'b0000000111100110;
            15'd3060: log10_cal = 16'b0000000111100110;
            15'd3061: log10_cal = 16'b0000000111100110;
            15'd3062: log10_cal = 16'b0000000111100111;
            15'd3063: log10_cal = 16'b0000000111100111;
            15'd3064: log10_cal = 16'b0000000111100111;
            15'd3065: log10_cal = 16'b0000000111100111;
            15'd3066: log10_cal = 16'b0000000111100111;
            15'd3067: log10_cal = 16'b0000000111100111;
            15'd3068: log10_cal = 16'b0000000111100111;
            15'd3069: log10_cal = 16'b0000000111101000;
            15'd3070: log10_cal = 16'b0000000111101000;
            15'd3071: log10_cal = 16'b0000000111101000;
            15'd3072: log10_cal = 16'b0000000111101000;
            15'd3073: log10_cal = 16'b0000000111101000;
            15'd3074: log10_cal = 16'b0000000111101000;
            15'd3075: log10_cal = 16'b0000000111101001;
            15'd3076: log10_cal = 16'b0000000111101001;
            15'd3077: log10_cal = 16'b0000000111101001;
            15'd3078: log10_cal = 16'b0000000111101001;
            15'd3079: log10_cal = 16'b0000000111101001;
            15'd3080: log10_cal = 16'b0000000111101001;
            15'd3081: log10_cal = 16'b0000000111101001;
            15'd3082: log10_cal = 16'b0000000111101010;
            15'd3083: log10_cal = 16'b0000000111101010;
            15'd3084: log10_cal = 16'b0000000111101010;
            15'd3085: log10_cal = 16'b0000000111101010;
            15'd3086: log10_cal = 16'b0000000111101010;
            15'd3087: log10_cal = 16'b0000000111101010;
            15'd3088: log10_cal = 16'b0000000111101010;
            15'd3089: log10_cal = 16'b0000000111101011;
            15'd3090: log10_cal = 16'b0000000111101011;
            15'd3091: log10_cal = 16'b0000000111101011;
            15'd3092: log10_cal = 16'b0000000111101011;
            15'd3093: log10_cal = 16'b0000000111101011;
            15'd3094: log10_cal = 16'b0000000111101011;
            15'd3095: log10_cal = 16'b0000000111101011;
            15'd3096: log10_cal = 16'b0000000111101100;
            15'd3097: log10_cal = 16'b0000000111101100;
            15'd3098: log10_cal = 16'b0000000111101100;
            15'd3099: log10_cal = 16'b0000000111101100;
            15'd3100: log10_cal = 16'b0000000111101100;
            15'd3101: log10_cal = 16'b0000000111101100;
            15'd3102: log10_cal = 16'b0000000111101100;
            15'd3103: log10_cal = 16'b0000000111101101;
            15'd3104: log10_cal = 16'b0000000111101101;
            15'd3105: log10_cal = 16'b0000000111101101;
            15'd3106: log10_cal = 16'b0000000111101101;
            15'd3107: log10_cal = 16'b0000000111101101;
            15'd3108: log10_cal = 16'b0000000111101101;
            15'd3109: log10_cal = 16'b0000000111101101;
            15'd3110: log10_cal = 16'b0000000111101110;
            15'd3111: log10_cal = 16'b0000000111101110;
            15'd3112: log10_cal = 16'b0000000111101110;
            15'd3113: log10_cal = 16'b0000000111101110;
            15'd3114: log10_cal = 16'b0000000111101110;
            15'd3115: log10_cal = 16'b0000000111101110;
            15'd3116: log10_cal = 16'b0000000111101110;
            15'd3117: log10_cal = 16'b0000000111101111;
            15'd3118: log10_cal = 16'b0000000111101111;
            15'd3119: log10_cal = 16'b0000000111101111;
            15'd3120: log10_cal = 16'b0000000111101111;
            15'd3121: log10_cal = 16'b0000000111101111;
            15'd3122: log10_cal = 16'b0000000111101111;
            15'd3123: log10_cal = 16'b0000000111101111;
            15'd3124: log10_cal = 16'b0000000111110000;
            15'd3125: log10_cal = 16'b0000000111110000;
            15'd3126: log10_cal = 16'b0000000111110000;
            15'd3127: log10_cal = 16'b0000000111110000;
            15'd3128: log10_cal = 16'b0000000111110000;
            15'd3129: log10_cal = 16'b0000000111110000;
            15'd3130: log10_cal = 16'b0000000111110000;
            15'd3131: log10_cal = 16'b0000000111110001;
            15'd3132: log10_cal = 16'b0000000111110001;
            15'd3133: log10_cal = 16'b0000000111110001;
            15'd3134: log10_cal = 16'b0000000111110001;
            15'd3135: log10_cal = 16'b0000000111110001;
            15'd3136: log10_cal = 16'b0000000111110001;
            15'd3137: log10_cal = 16'b0000000111110001;
            15'd3138: log10_cal = 16'b0000000111110010;
            15'd3139: log10_cal = 16'b0000000111110010;
            15'd3140: log10_cal = 16'b0000000111110010;
            15'd3141: log10_cal = 16'b0000000111110010;
            15'd3142: log10_cal = 16'b0000000111110010;
            15'd3143: log10_cal = 16'b0000000111110010;
            15'd3144: log10_cal = 16'b0000000111110010;
            15'd3145: log10_cal = 16'b0000000111110011;
            15'd3146: log10_cal = 16'b0000000111110011;
            15'd3147: log10_cal = 16'b0000000111110011;
            15'd3148: log10_cal = 16'b0000000111110011;
            15'd3149: log10_cal = 16'b0000000111110011;
            15'd3150: log10_cal = 16'b0000000111110011;
            15'd3151: log10_cal = 16'b0000000111110011;
            15'd3152: log10_cal = 16'b0000000111110100;
            15'd3153: log10_cal = 16'b0000000111110100;
            15'd3154: log10_cal = 16'b0000000111110100;
            15'd3155: log10_cal = 16'b0000000111110100;
            15'd3156: log10_cal = 16'b0000000111110100;
            15'd3157: log10_cal = 16'b0000000111110100;
            15'd3158: log10_cal = 16'b0000000111110100;
            15'd3159: log10_cal = 16'b0000000111110100;
            15'd3160: log10_cal = 16'b0000000111110101;
            15'd3161: log10_cal = 16'b0000000111110101;
            15'd3162: log10_cal = 16'b0000000111110101;
            15'd3163: log10_cal = 16'b0000000111110101;
            15'd3164: log10_cal = 16'b0000000111110101;
            15'd3165: log10_cal = 16'b0000000111110101;
            15'd3166: log10_cal = 16'b0000000111110101;
            15'd3167: log10_cal = 16'b0000000111110110;
            15'd3168: log10_cal = 16'b0000000111110110;
            15'd3169: log10_cal = 16'b0000000111110110;
            15'd3170: log10_cal = 16'b0000000111110110;
            15'd3171: log10_cal = 16'b0000000111110110;
            15'd3172: log10_cal = 16'b0000000111110110;
            15'd3173: log10_cal = 16'b0000000111110110;
            15'd3174: log10_cal = 16'b0000000111110111;
            15'd3175: log10_cal = 16'b0000000111110111;
            15'd3176: log10_cal = 16'b0000000111110111;
            15'd3177: log10_cal = 16'b0000000111110111;
            15'd3178: log10_cal = 16'b0000000111110111;
            15'd3179: log10_cal = 16'b0000000111110111;
            15'd3180: log10_cal = 16'b0000000111110111;
            15'd3181: log10_cal = 16'b0000000111111000;
            15'd3182: log10_cal = 16'b0000000111111000;
            15'd3183: log10_cal = 16'b0000000111111000;
            15'd3184: log10_cal = 16'b0000000111111000;
            15'd3185: log10_cal = 16'b0000000111111000;
            15'd3186: log10_cal = 16'b0000000111111000;
            15'd3187: log10_cal = 16'b0000000111111000;
            15'd3188: log10_cal = 16'b0000000111111001;
            15'd3189: log10_cal = 16'b0000000111111001;
            15'd3190: log10_cal = 16'b0000000111111001;
            15'd3191: log10_cal = 16'b0000000111111001;
            15'd3192: log10_cal = 16'b0000000111111001;
            15'd3193: log10_cal = 16'b0000000111111001;
            15'd3194: log10_cal = 16'b0000000111111001;
            15'd3195: log10_cal = 16'b0000000111111010;
            15'd3196: log10_cal = 16'b0000000111111010;
            15'd3197: log10_cal = 16'b0000000111111010;
            15'd3198: log10_cal = 16'b0000000111111010;
            15'd3199: log10_cal = 16'b0000000111111010;
            15'd3200: log10_cal = 16'b0000000111111010;
            15'd3201: log10_cal = 16'b0000000111111010;
            15'd3202: log10_cal = 16'b0000000111111011;
            15'd3203: log10_cal = 16'b0000000111111011;
            15'd3204: log10_cal = 16'b0000000111111011;
            15'd3205: log10_cal = 16'b0000000111111011;
            15'd3206: log10_cal = 16'b0000000111111011;
            15'd3207: log10_cal = 16'b0000000111111011;
            15'd3208: log10_cal = 16'b0000000111111011;
            15'd3209: log10_cal = 16'b0000000111111011;
            15'd3210: log10_cal = 16'b0000000111111100;
            15'd3211: log10_cal = 16'b0000000111111100;
            15'd3212: log10_cal = 16'b0000000111111100;
            15'd3213: log10_cal = 16'b0000000111111100;
            15'd3214: log10_cal = 16'b0000000111111100;
            15'd3215: log10_cal = 16'b0000000111111100;
            15'd3216: log10_cal = 16'b0000000111111100;
            15'd3217: log10_cal = 16'b0000000111111101;
            15'd3218: log10_cal = 16'b0000000111111101;
            15'd3219: log10_cal = 16'b0000000111111101;
            15'd3220: log10_cal = 16'b0000000111111101;
            15'd3221: log10_cal = 16'b0000000111111101;
            15'd3222: log10_cal = 16'b0000000111111101;
            15'd3223: log10_cal = 16'b0000000111111101;
            15'd3224: log10_cal = 16'b0000000111111110;
            15'd3225: log10_cal = 16'b0000000111111110;
            15'd3226: log10_cal = 16'b0000000111111110;
            15'd3227: log10_cal = 16'b0000000111111110;
            15'd3228: log10_cal = 16'b0000000111111110;
            15'd3229: log10_cal = 16'b0000000111111110;
            15'd3230: log10_cal = 16'b0000000111111110;
            15'd3231: log10_cal = 16'b0000000111111111;
            15'd3232: log10_cal = 16'b0000000111111111;
            15'd3233: log10_cal = 16'b0000000111111111;
            15'd3234: log10_cal = 16'b0000000111111111;
            15'd3235: log10_cal = 16'b0000000111111111;
            15'd3236: log10_cal = 16'b0000000111111111;
            15'd3237: log10_cal = 16'b0000000111111111;
            15'd3238: log10_cal = 16'b0000000111111111;
            15'd3239: log10_cal = 16'b0000001000000000;
            15'd3240: log10_cal = 16'b0000001000000000;
            15'd3241: log10_cal = 16'b0000001000000000;
            15'd3242: log10_cal = 16'b0000001000000000;
            15'd3243: log10_cal = 16'b0000001000000000;
            15'd3244: log10_cal = 16'b0000001000000000;
            15'd3245: log10_cal = 16'b0000001000000000;
            15'd3246: log10_cal = 16'b0000001000000001;
            15'd3247: log10_cal = 16'b0000001000000001;
            15'd3248: log10_cal = 16'b0000001000000001;
            15'd3249: log10_cal = 16'b0000001000000001;
            15'd3250: log10_cal = 16'b0000001000000001;
            15'd3251: log10_cal = 16'b0000001000000001;
            15'd3252: log10_cal = 16'b0000001000000001;
            15'd3253: log10_cal = 16'b0000001000000010;
            15'd3254: log10_cal = 16'b0000001000000010;
            15'd3255: log10_cal = 16'b0000001000000010;
            15'd3256: log10_cal = 16'b0000001000000010;
            15'd3257: log10_cal = 16'b0000001000000010;
            15'd3258: log10_cal = 16'b0000001000000010;
            15'd3259: log10_cal = 16'b0000001000000010;
            15'd3260: log10_cal = 16'b0000001000000010;
            15'd3261: log10_cal = 16'b0000001000000011;
            15'd3262: log10_cal = 16'b0000001000000011;
            15'd3263: log10_cal = 16'b0000001000000011;
            15'd3264: log10_cal = 16'b0000001000000011;
            15'd3265: log10_cal = 16'b0000001000000011;
            15'd3266: log10_cal = 16'b0000001000000011;
            15'd3267: log10_cal = 16'b0000001000000011;
            15'd3268: log10_cal = 16'b0000001000000100;
            15'd3269: log10_cal = 16'b0000001000000100;
            15'd3270: log10_cal = 16'b0000001000000100;
            15'd3271: log10_cal = 16'b0000001000000100;
            15'd3272: log10_cal = 16'b0000001000000100;
            15'd3273: log10_cal = 16'b0000001000000100;
            15'd3274: log10_cal = 16'b0000001000000100;
            15'd3275: log10_cal = 16'b0000001000000101;
            15'd3276: log10_cal = 16'b0000001000000101;
            15'd3277: log10_cal = 16'b0000001000000101;
            15'd3278: log10_cal = 16'b0000001000000101;
            15'd3279: log10_cal = 16'b0000001000000101;
            15'd3280: log10_cal = 16'b0000001000000101;
            15'd3281: log10_cal = 16'b0000001000000101;
            15'd3282: log10_cal = 16'b0000001000000101;
            15'd3283: log10_cal = 16'b0000001000000110;
            15'd3284: log10_cal = 16'b0000001000000110;
            15'd3285: log10_cal = 16'b0000001000000110;
            15'd3286: log10_cal = 16'b0000001000000110;
            15'd3287: log10_cal = 16'b0000001000000110;
            15'd3288: log10_cal = 16'b0000001000000110;
            15'd3289: log10_cal = 16'b0000001000000110;
            15'd3290: log10_cal = 16'b0000001000000111;
            15'd3291: log10_cal = 16'b0000001000000111;
            15'd3292: log10_cal = 16'b0000001000000111;
            15'd3293: log10_cal = 16'b0000001000000111;
            15'd3294: log10_cal = 16'b0000001000000111;
            15'd3295: log10_cal = 16'b0000001000000111;
            15'd3296: log10_cal = 16'b0000001000000111;
            15'd3297: log10_cal = 16'b0000001000001000;
            15'd3298: log10_cal = 16'b0000001000001000;
            15'd3299: log10_cal = 16'b0000001000001000;
            15'd3300: log10_cal = 16'b0000001000001000;
            15'd3301: log10_cal = 16'b0000001000001000;
            15'd3302: log10_cal = 16'b0000001000001000;
            15'd3303: log10_cal = 16'b0000001000001000;
            15'd3304: log10_cal = 16'b0000001000001000;
            15'd3305: log10_cal = 16'b0000001000001001;
            15'd3306: log10_cal = 16'b0000001000001001;
            15'd3307: log10_cal = 16'b0000001000001001;
            15'd3308: log10_cal = 16'b0000001000001001;
            15'd3309: log10_cal = 16'b0000001000001001;
            15'd3310: log10_cal = 16'b0000001000001001;
            15'd3311: log10_cal = 16'b0000001000001001;
            15'd3312: log10_cal = 16'b0000001000001010;
            15'd3313: log10_cal = 16'b0000001000001010;
            15'd3314: log10_cal = 16'b0000001000001010;
            15'd3315: log10_cal = 16'b0000001000001010;
            15'd3316: log10_cal = 16'b0000001000001010;
            15'd3317: log10_cal = 16'b0000001000001010;
            15'd3318: log10_cal = 16'b0000001000001010;
            15'd3319: log10_cal = 16'b0000001000001010;
            15'd3320: log10_cal = 16'b0000001000001011;
            15'd3321: log10_cal = 16'b0000001000001011;
            15'd3322: log10_cal = 16'b0000001000001011;
            15'd3323: log10_cal = 16'b0000001000001011;
            15'd3324: log10_cal = 16'b0000001000001011;
            15'd3325: log10_cal = 16'b0000001000001011;
            15'd3326: log10_cal = 16'b0000001000001011;
            15'd3327: log10_cal = 16'b0000001000001100;
            15'd3328: log10_cal = 16'b0000001000001100;
            15'd3329: log10_cal = 16'b0000001000001100;
            15'd3330: log10_cal = 16'b0000001000001100;
            15'd3331: log10_cal = 16'b0000001000001100;
            15'd3332: log10_cal = 16'b0000001000001100;
            15'd3333: log10_cal = 16'b0000001000001100;
            15'd3334: log10_cal = 16'b0000001000001100;
            15'd3335: log10_cal = 16'b0000001000001101;
            15'd3336: log10_cal = 16'b0000001000001101;
            15'd3337: log10_cal = 16'b0000001000001101;
            15'd3338: log10_cal = 16'b0000001000001101;
            15'd3339: log10_cal = 16'b0000001000001101;
            15'd3340: log10_cal = 16'b0000001000001101;
            15'd3341: log10_cal = 16'b0000001000001101;
            15'd3342: log10_cal = 16'b0000001000001110;
            15'd3343: log10_cal = 16'b0000001000001110;
            15'd3344: log10_cal = 16'b0000001000001110;
            15'd3345: log10_cal = 16'b0000001000001110;
            15'd3346: log10_cal = 16'b0000001000001110;
            15'd3347: log10_cal = 16'b0000001000001110;
            15'd3348: log10_cal = 16'b0000001000001110;
            15'd3349: log10_cal = 16'b0000001000001110;
            15'd3350: log10_cal = 16'b0000001000001111;
            15'd3351: log10_cal = 16'b0000001000001111;
            15'd3352: log10_cal = 16'b0000001000001111;
            15'd3353: log10_cal = 16'b0000001000001111;
            15'd3354: log10_cal = 16'b0000001000001111;
            15'd3355: log10_cal = 16'b0000001000001111;
            15'd3356: log10_cal = 16'b0000001000001111;
            15'd3357: log10_cal = 16'b0000001000010000;
            15'd3358: log10_cal = 16'b0000001000010000;
            15'd3359: log10_cal = 16'b0000001000010000;
            15'd3360: log10_cal = 16'b0000001000010000;
            15'd3361: log10_cal = 16'b0000001000010000;
            15'd3362: log10_cal = 16'b0000001000010000;
            15'd3363: log10_cal = 16'b0000001000010000;
            15'd3364: log10_cal = 16'b0000001000010000;
            15'd3365: log10_cal = 16'b0000001000010001;
            15'd3366: log10_cal = 16'b0000001000010001;
            15'd3367: log10_cal = 16'b0000001000010001;
            15'd3368: log10_cal = 16'b0000001000010001;
            15'd3369: log10_cal = 16'b0000001000010001;
            15'd3370: log10_cal = 16'b0000001000010001;
            15'd3371: log10_cal = 16'b0000001000010001;
            15'd3372: log10_cal = 16'b0000001000010010;
            15'd3373: log10_cal = 16'b0000001000010010;
            15'd3374: log10_cal = 16'b0000001000010010;
            15'd3375: log10_cal = 16'b0000001000010010;
            15'd3376: log10_cal = 16'b0000001000010010;
            15'd3377: log10_cal = 16'b0000001000010010;
            15'd3378: log10_cal = 16'b0000001000010010;
            15'd3379: log10_cal = 16'b0000001000010010;
            15'd3380: log10_cal = 16'b0000001000010011;
            15'd3381: log10_cal = 16'b0000001000010011;
            15'd3382: log10_cal = 16'b0000001000010011;
            15'd3383: log10_cal = 16'b0000001000010011;
            15'd3384: log10_cal = 16'b0000001000010011;
            15'd3385: log10_cal = 16'b0000001000010011;
            15'd3386: log10_cal = 16'b0000001000010011;
            15'd3387: log10_cal = 16'b0000001000010011;
            15'd3388: log10_cal = 16'b0000001000010100;
            15'd3389: log10_cal = 16'b0000001000010100;
            15'd3390: log10_cal = 16'b0000001000010100;
            15'd3391: log10_cal = 16'b0000001000010100;
            15'd3392: log10_cal = 16'b0000001000010100;
            15'd3393: log10_cal = 16'b0000001000010100;
            15'd3394: log10_cal = 16'b0000001000010100;
            15'd3395: log10_cal = 16'b0000001000010101;
            15'd3396: log10_cal = 16'b0000001000010101;
            15'd3397: log10_cal = 16'b0000001000010101;
            15'd3398: log10_cal = 16'b0000001000010101;
            15'd3399: log10_cal = 16'b0000001000010101;
            15'd3400: log10_cal = 16'b0000001000010101;
            15'd3401: log10_cal = 16'b0000001000010101;
            15'd3402: log10_cal = 16'b0000001000010101;
            15'd3403: log10_cal = 16'b0000001000010110;
            15'd3404: log10_cal = 16'b0000001000010110;
            15'd3405: log10_cal = 16'b0000001000010110;
            15'd3406: log10_cal = 16'b0000001000010110;
            15'd3407: log10_cal = 16'b0000001000010110;
            15'd3408: log10_cal = 16'b0000001000010110;
            15'd3409: log10_cal = 16'b0000001000010110;
            15'd3410: log10_cal = 16'b0000001000010110;
            15'd3411: log10_cal = 16'b0000001000010111;
            15'd3412: log10_cal = 16'b0000001000010111;
            15'd3413: log10_cal = 16'b0000001000010111;
            15'd3414: log10_cal = 16'b0000001000010111;
            15'd3415: log10_cal = 16'b0000001000010111;
            15'd3416: log10_cal = 16'b0000001000010111;
            15'd3417: log10_cal = 16'b0000001000010111;
            15'd3418: log10_cal = 16'b0000001000011000;
            15'd3419: log10_cal = 16'b0000001000011000;
            15'd3420: log10_cal = 16'b0000001000011000;
            15'd3421: log10_cal = 16'b0000001000011000;
            15'd3422: log10_cal = 16'b0000001000011000;
            15'd3423: log10_cal = 16'b0000001000011000;
            15'd3424: log10_cal = 16'b0000001000011000;
            15'd3425: log10_cal = 16'b0000001000011000;
            15'd3426: log10_cal = 16'b0000001000011001;
            15'd3427: log10_cal = 16'b0000001000011001;
            15'd3428: log10_cal = 16'b0000001000011001;
            15'd3429: log10_cal = 16'b0000001000011001;
            15'd3430: log10_cal = 16'b0000001000011001;
            15'd3431: log10_cal = 16'b0000001000011001;
            15'd3432: log10_cal = 16'b0000001000011001;
            15'd3433: log10_cal = 16'b0000001000011001;
            15'd3434: log10_cal = 16'b0000001000011010;
            15'd3435: log10_cal = 16'b0000001000011010;
            15'd3436: log10_cal = 16'b0000001000011010;
            15'd3437: log10_cal = 16'b0000001000011010;
            15'd3438: log10_cal = 16'b0000001000011010;
            15'd3439: log10_cal = 16'b0000001000011010;
            15'd3440: log10_cal = 16'b0000001000011010;
            15'd3441: log10_cal = 16'b0000001000011011;
            15'd3442: log10_cal = 16'b0000001000011011;
            15'd3443: log10_cal = 16'b0000001000011011;
            15'd3444: log10_cal = 16'b0000001000011011;
            15'd3445: log10_cal = 16'b0000001000011011;
            15'd3446: log10_cal = 16'b0000001000011011;
            15'd3447: log10_cal = 16'b0000001000011011;
            15'd3448: log10_cal = 16'b0000001000011011;
            15'd3449: log10_cal = 16'b0000001000011100;
            15'd3450: log10_cal = 16'b0000001000011100;
            15'd3451: log10_cal = 16'b0000001000011100;
            15'd3452: log10_cal = 16'b0000001000011100;
            15'd3453: log10_cal = 16'b0000001000011100;
            15'd3454: log10_cal = 16'b0000001000011100;
            15'd3455: log10_cal = 16'b0000001000011100;
            15'd3456: log10_cal = 16'b0000001000011100;
            15'd3457: log10_cal = 16'b0000001000011101;
            15'd3458: log10_cal = 16'b0000001000011101;
            15'd3459: log10_cal = 16'b0000001000011101;
            15'd3460: log10_cal = 16'b0000001000011101;
            15'd3461: log10_cal = 16'b0000001000011101;
            15'd3462: log10_cal = 16'b0000001000011101;
            15'd3463: log10_cal = 16'b0000001000011101;
            15'd3464: log10_cal = 16'b0000001000011101;
            15'd3465: log10_cal = 16'b0000001000011110;
            15'd3466: log10_cal = 16'b0000001000011110;
            15'd3467: log10_cal = 16'b0000001000011110;
            15'd3468: log10_cal = 16'b0000001000011110;
            15'd3469: log10_cal = 16'b0000001000011110;
            15'd3470: log10_cal = 16'b0000001000011110;
            15'd3471: log10_cal = 16'b0000001000011110;
            15'd3472: log10_cal = 16'b0000001000011111;
            15'd3473: log10_cal = 16'b0000001000011111;
            15'd3474: log10_cal = 16'b0000001000011111;
            15'd3475: log10_cal = 16'b0000001000011111;
            15'd3476: log10_cal = 16'b0000001000011111;
            15'd3477: log10_cal = 16'b0000001000011111;
            15'd3478: log10_cal = 16'b0000001000011111;
            15'd3479: log10_cal = 16'b0000001000011111;
            15'd3480: log10_cal = 16'b0000001000100000;
            15'd3481: log10_cal = 16'b0000001000100000;
            15'd3482: log10_cal = 16'b0000001000100000;
            15'd3483: log10_cal = 16'b0000001000100000;
            15'd3484: log10_cal = 16'b0000001000100000;
            15'd3485: log10_cal = 16'b0000001000100000;
            15'd3486: log10_cal = 16'b0000001000100000;
            15'd3487: log10_cal = 16'b0000001000100000;
            15'd3488: log10_cal = 16'b0000001000100001;
            15'd3489: log10_cal = 16'b0000001000100001;
            15'd3490: log10_cal = 16'b0000001000100001;
            15'd3491: log10_cal = 16'b0000001000100001;
            15'd3492: log10_cal = 16'b0000001000100001;
            15'd3493: log10_cal = 16'b0000001000100001;
            15'd3494: log10_cal = 16'b0000001000100001;
            15'd3495: log10_cal = 16'b0000001000100001;
            15'd3496: log10_cal = 16'b0000001000100010;
            15'd3497: log10_cal = 16'b0000001000100010;
            15'd3498: log10_cal = 16'b0000001000100010;
            15'd3499: log10_cal = 16'b0000001000100010;
            15'd3500: log10_cal = 16'b0000001000100010;
            15'd3501: log10_cal = 16'b0000001000100010;
            15'd3502: log10_cal = 16'b0000001000100010;
            15'd3503: log10_cal = 16'b0000001000100010;
            15'd3504: log10_cal = 16'b0000001000100011;
            15'd3505: log10_cal = 16'b0000001000100011;
            15'd3506: log10_cal = 16'b0000001000100011;
            15'd3507: log10_cal = 16'b0000001000100011;
            15'd3508: log10_cal = 16'b0000001000100011;
            15'd3509: log10_cal = 16'b0000001000100011;
            15'd3510: log10_cal = 16'b0000001000100011;
            15'd3511: log10_cal = 16'b0000001000100011;
            15'd3512: log10_cal = 16'b0000001000100100;
            15'd3513: log10_cal = 16'b0000001000100100;
            15'd3514: log10_cal = 16'b0000001000100100;
            15'd3515: log10_cal = 16'b0000001000100100;
            15'd3516: log10_cal = 16'b0000001000100100;
            15'd3517: log10_cal = 16'b0000001000100100;
            15'd3518: log10_cal = 16'b0000001000100100;
            15'd3519: log10_cal = 16'b0000001000100100;
            15'd3520: log10_cal = 16'b0000001000100101;
            15'd3521: log10_cal = 16'b0000001000100101;
            15'd3522: log10_cal = 16'b0000001000100101;
            15'd3523: log10_cal = 16'b0000001000100101;
            15'd3524: log10_cal = 16'b0000001000100101;
            15'd3525: log10_cal = 16'b0000001000100101;
            15'd3526: log10_cal = 16'b0000001000100101;
            15'd3527: log10_cal = 16'b0000001000100101;
            15'd3528: log10_cal = 16'b0000001000100110;
            15'd3529: log10_cal = 16'b0000001000100110;
            15'd3530: log10_cal = 16'b0000001000100110;
            15'd3531: log10_cal = 16'b0000001000100110;
            15'd3532: log10_cal = 16'b0000001000100110;
            15'd3533: log10_cal = 16'b0000001000100110;
            15'd3534: log10_cal = 16'b0000001000100110;
            15'd3535: log10_cal = 16'b0000001000100111;
            15'd3536: log10_cal = 16'b0000001000100111;
            15'd3537: log10_cal = 16'b0000001000100111;
            15'd3538: log10_cal = 16'b0000001000100111;
            15'd3539: log10_cal = 16'b0000001000100111;
            15'd3540: log10_cal = 16'b0000001000100111;
            15'd3541: log10_cal = 16'b0000001000100111;
            15'd3542: log10_cal = 16'b0000001000100111;
            15'd3543: log10_cal = 16'b0000001000101000;
            15'd3544: log10_cal = 16'b0000001000101000;
            15'd3545: log10_cal = 16'b0000001000101000;
            15'd3546: log10_cal = 16'b0000001000101000;
            15'd3547: log10_cal = 16'b0000001000101000;
            15'd3548: log10_cal = 16'b0000001000101000;
            15'd3549: log10_cal = 16'b0000001000101000;
            15'd3550: log10_cal = 16'b0000001000101000;
            15'd3551: log10_cal = 16'b0000001000101001;
            15'd3552: log10_cal = 16'b0000001000101001;
            15'd3553: log10_cal = 16'b0000001000101001;
            15'd3554: log10_cal = 16'b0000001000101001;
            15'd3555: log10_cal = 16'b0000001000101001;
            15'd3556: log10_cal = 16'b0000001000101001;
            15'd3557: log10_cal = 16'b0000001000101001;
            15'd3558: log10_cal = 16'b0000001000101001;
            15'd3559: log10_cal = 16'b0000001000101010;
            15'd3560: log10_cal = 16'b0000001000101010;
            15'd3561: log10_cal = 16'b0000001000101010;
            15'd3562: log10_cal = 16'b0000001000101010;
            15'd3563: log10_cal = 16'b0000001000101010;
            15'd3564: log10_cal = 16'b0000001000101010;
            15'd3565: log10_cal = 16'b0000001000101010;
            15'd3566: log10_cal = 16'b0000001000101010;
            15'd3567: log10_cal = 16'b0000001000101011;
            15'd3568: log10_cal = 16'b0000001000101011;
            15'd3569: log10_cal = 16'b0000001000101011;
            15'd3570: log10_cal = 16'b0000001000101011;
            15'd3571: log10_cal = 16'b0000001000101011;
            15'd3572: log10_cal = 16'b0000001000101011;
            15'd3573: log10_cal = 16'b0000001000101011;
            15'd3574: log10_cal = 16'b0000001000101011;
            15'd3575: log10_cal = 16'b0000001000101100;
            15'd3576: log10_cal = 16'b0000001000101100;
            15'd3577: log10_cal = 16'b0000001000101100;
            15'd3578: log10_cal = 16'b0000001000101100;
            15'd3579: log10_cal = 16'b0000001000101100;
            15'd3580: log10_cal = 16'b0000001000101100;
            15'd3581: log10_cal = 16'b0000001000101100;
            15'd3582: log10_cal = 16'b0000001000101100;
            15'd3583: log10_cal = 16'b0000001000101101;
            15'd3584: log10_cal = 16'b0000001000101101;
            15'd3585: log10_cal = 16'b0000001000101101;
            15'd3586: log10_cal = 16'b0000001000101101;
            15'd3587: log10_cal = 16'b0000001000101101;
            15'd3588: log10_cal = 16'b0000001000101101;
            15'd3589: log10_cal = 16'b0000001000101101;
            15'd3590: log10_cal = 16'b0000001000101101;
            15'd3591: log10_cal = 16'b0000001000101101;
            15'd3592: log10_cal = 16'b0000001000101110;
            15'd3593: log10_cal = 16'b0000001000101110;
            15'd3594: log10_cal = 16'b0000001000101110;
            15'd3595: log10_cal = 16'b0000001000101110;
            15'd3596: log10_cal = 16'b0000001000101110;
            15'd3597: log10_cal = 16'b0000001000101110;
            15'd3598: log10_cal = 16'b0000001000101110;
            15'd3599: log10_cal = 16'b0000001000101110;
            15'd3600: log10_cal = 16'b0000001000101111;
            15'd3601: log10_cal = 16'b0000001000101111;
            15'd3602: log10_cal = 16'b0000001000101111;
            15'd3603: log10_cal = 16'b0000001000101111;
            15'd3604: log10_cal = 16'b0000001000101111;
            15'd3605: log10_cal = 16'b0000001000101111;
            15'd3606: log10_cal = 16'b0000001000101111;
            15'd3607: log10_cal = 16'b0000001000101111;
            15'd3608: log10_cal = 16'b0000001000110000;
            15'd3609: log10_cal = 16'b0000001000110000;
            15'd3610: log10_cal = 16'b0000001000110000;
            15'd3611: log10_cal = 16'b0000001000110000;
            15'd3612: log10_cal = 16'b0000001000110000;
            15'd3613: log10_cal = 16'b0000001000110000;
            15'd3614: log10_cal = 16'b0000001000110000;
            15'd3615: log10_cal = 16'b0000001000110000;
            15'd3616: log10_cal = 16'b0000001000110001;
            15'd3617: log10_cal = 16'b0000001000110001;
            15'd3618: log10_cal = 16'b0000001000110001;
            15'd3619: log10_cal = 16'b0000001000110001;
            15'd3620: log10_cal = 16'b0000001000110001;
            15'd3621: log10_cal = 16'b0000001000110001;
            15'd3622: log10_cal = 16'b0000001000110001;
            15'd3623: log10_cal = 16'b0000001000110001;
            15'd3624: log10_cal = 16'b0000001000110010;
            15'd3625: log10_cal = 16'b0000001000110010;
            15'd3626: log10_cal = 16'b0000001000110010;
            15'd3627: log10_cal = 16'b0000001000110010;
            15'd3628: log10_cal = 16'b0000001000110010;
            15'd3629: log10_cal = 16'b0000001000110010;
            15'd3630: log10_cal = 16'b0000001000110010;
            15'd3631: log10_cal = 16'b0000001000110010;
            15'd3632: log10_cal = 16'b0000001000110011;
            15'd3633: log10_cal = 16'b0000001000110011;
            15'd3634: log10_cal = 16'b0000001000110011;
            15'd3635: log10_cal = 16'b0000001000110011;
            15'd3636: log10_cal = 16'b0000001000110011;
            15'd3637: log10_cal = 16'b0000001000110011;
            15'd3638: log10_cal = 16'b0000001000110011;
            15'd3639: log10_cal = 16'b0000001000110011;
            15'd3640: log10_cal = 16'b0000001000110100;
            15'd3641: log10_cal = 16'b0000001000110100;
            15'd3642: log10_cal = 16'b0000001000110100;
            15'd3643: log10_cal = 16'b0000001000110100;
            15'd3644: log10_cal = 16'b0000001000110100;
            15'd3645: log10_cal = 16'b0000001000110100;
            15'd3646: log10_cal = 16'b0000001000110100;
            15'd3647: log10_cal = 16'b0000001000110100;
            15'd3648: log10_cal = 16'b0000001000110100;
            15'd3649: log10_cal = 16'b0000001000110101;
            15'd3650: log10_cal = 16'b0000001000110101;
            15'd3651: log10_cal = 16'b0000001000110101;
            15'd3652: log10_cal = 16'b0000001000110101;
            15'd3653: log10_cal = 16'b0000001000110101;
            15'd3654: log10_cal = 16'b0000001000110101;
            15'd3655: log10_cal = 16'b0000001000110101;
            15'd3656: log10_cal = 16'b0000001000110101;
            15'd3657: log10_cal = 16'b0000001000110110;
            15'd3658: log10_cal = 16'b0000001000110110;
            15'd3659: log10_cal = 16'b0000001000110110;
            15'd3660: log10_cal = 16'b0000001000110110;
            15'd3661: log10_cal = 16'b0000001000110110;
            15'd3662: log10_cal = 16'b0000001000110110;
            15'd3663: log10_cal = 16'b0000001000110110;
            15'd3664: log10_cal = 16'b0000001000110110;
            15'd3665: log10_cal = 16'b0000001000110111;
            15'd3666: log10_cal = 16'b0000001000110111;
            15'd3667: log10_cal = 16'b0000001000110111;
            15'd3668: log10_cal = 16'b0000001000110111;
            15'd3669: log10_cal = 16'b0000001000110111;
            15'd3670: log10_cal = 16'b0000001000110111;
            15'd3671: log10_cal = 16'b0000001000110111;
            15'd3672: log10_cal = 16'b0000001000110111;
            15'd3673: log10_cal = 16'b0000001000111000;
            15'd3674: log10_cal = 16'b0000001000111000;
            15'd3675: log10_cal = 16'b0000001000111000;
            15'd3676: log10_cal = 16'b0000001000111000;
            15'd3677: log10_cal = 16'b0000001000111000;
            15'd3678: log10_cal = 16'b0000001000111000;
            15'd3679: log10_cal = 16'b0000001000111000;
            15'd3680: log10_cal = 16'b0000001000111000;
            15'd3681: log10_cal = 16'b0000001000111001;
            15'd3682: log10_cal = 16'b0000001000111001;
            15'd3683: log10_cal = 16'b0000001000111001;
            15'd3684: log10_cal = 16'b0000001000111001;
            15'd3685: log10_cal = 16'b0000001000111001;
            15'd3686: log10_cal = 16'b0000001000111001;
            15'd3687: log10_cal = 16'b0000001000111001;
            15'd3688: log10_cal = 16'b0000001000111001;
            15'd3689: log10_cal = 16'b0000001000111001;
            15'd3690: log10_cal = 16'b0000001000111010;
            15'd3691: log10_cal = 16'b0000001000111010;
            15'd3692: log10_cal = 16'b0000001000111010;
            15'd3693: log10_cal = 16'b0000001000111010;
            15'd3694: log10_cal = 16'b0000001000111010;
            15'd3695: log10_cal = 16'b0000001000111010;
            15'd3696: log10_cal = 16'b0000001000111010;
            15'd3697: log10_cal = 16'b0000001000111010;
            15'd3698: log10_cal = 16'b0000001000111011;
            15'd3699: log10_cal = 16'b0000001000111011;
            15'd3700: log10_cal = 16'b0000001000111011;
            15'd3701: log10_cal = 16'b0000001000111011;
            15'd3702: log10_cal = 16'b0000001000111011;
            15'd3703: log10_cal = 16'b0000001000111011;
            15'd3704: log10_cal = 16'b0000001000111011;
            15'd3705: log10_cal = 16'b0000001000111011;
            15'd3706: log10_cal = 16'b0000001000111100;
            15'd3707: log10_cal = 16'b0000001000111100;
            15'd3708: log10_cal = 16'b0000001000111100;
            15'd3709: log10_cal = 16'b0000001000111100;
            15'd3710: log10_cal = 16'b0000001000111100;
            15'd3711: log10_cal = 16'b0000001000111100;
            15'd3712: log10_cal = 16'b0000001000111100;
            15'd3713: log10_cal = 16'b0000001000111100;
            15'd3714: log10_cal = 16'b0000001000111100;
            15'd3715: log10_cal = 16'b0000001000111101;
            15'd3716: log10_cal = 16'b0000001000111101;
            15'd3717: log10_cal = 16'b0000001000111101;
            15'd3718: log10_cal = 16'b0000001000111101;
            15'd3719: log10_cal = 16'b0000001000111101;
            15'd3720: log10_cal = 16'b0000001000111101;
            15'd3721: log10_cal = 16'b0000001000111101;
            15'd3722: log10_cal = 16'b0000001000111101;
            15'd3723: log10_cal = 16'b0000001000111110;
            15'd3724: log10_cal = 16'b0000001000111110;
            15'd3725: log10_cal = 16'b0000001000111110;
            15'd3726: log10_cal = 16'b0000001000111110;
            15'd3727: log10_cal = 16'b0000001000111110;
            15'd3728: log10_cal = 16'b0000001000111110;
            15'd3729: log10_cal = 16'b0000001000111110;
            15'd3730: log10_cal = 16'b0000001000111110;
            15'd3731: log10_cal = 16'b0000001000111111;
            15'd3732: log10_cal = 16'b0000001000111111;
            15'd3733: log10_cal = 16'b0000001000111111;
            15'd3734: log10_cal = 16'b0000001000111111;
            15'd3735: log10_cal = 16'b0000001000111111;
            15'd3736: log10_cal = 16'b0000001000111111;
            15'd3737: log10_cal = 16'b0000001000111111;
            15'd3738: log10_cal = 16'b0000001000111111;
            15'd3739: log10_cal = 16'b0000001000111111;
            15'd3740: log10_cal = 16'b0000001001000000;
            15'd3741: log10_cal = 16'b0000001001000000;
            15'd3742: log10_cal = 16'b0000001001000000;
            15'd3743: log10_cal = 16'b0000001001000000;
            15'd3744: log10_cal = 16'b0000001001000000;
            15'd3745: log10_cal = 16'b0000001001000000;
            15'd3746: log10_cal = 16'b0000001001000000;
            15'd3747: log10_cal = 16'b0000001001000000;
            15'd3748: log10_cal = 16'b0000001001000001;
            15'd3749: log10_cal = 16'b0000001001000001;
            15'd3750: log10_cal = 16'b0000001001000001;
            15'd3751: log10_cal = 16'b0000001001000001;
            15'd3752: log10_cal = 16'b0000001001000001;
            15'd3753: log10_cal = 16'b0000001001000001;
            15'd3754: log10_cal = 16'b0000001001000001;
            15'd3755: log10_cal = 16'b0000001001000001;
            15'd3756: log10_cal = 16'b0000001001000001;
            15'd3757: log10_cal = 16'b0000001001000010;
            15'd3758: log10_cal = 16'b0000001001000010;
            15'd3759: log10_cal = 16'b0000001001000010;
            15'd3760: log10_cal = 16'b0000001001000010;
            15'd3761: log10_cal = 16'b0000001001000010;
            15'd3762: log10_cal = 16'b0000001001000010;
            15'd3763: log10_cal = 16'b0000001001000010;
            15'd3764: log10_cal = 16'b0000001001000010;
            15'd3765: log10_cal = 16'b0000001001000011;
            15'd3766: log10_cal = 16'b0000001001000011;
            15'd3767: log10_cal = 16'b0000001001000011;
            15'd3768: log10_cal = 16'b0000001001000011;
            15'd3769: log10_cal = 16'b0000001001000011;
            15'd3770: log10_cal = 16'b0000001001000011;
            15'd3771: log10_cal = 16'b0000001001000011;
            15'd3772: log10_cal = 16'b0000001001000011;
            15'd3773: log10_cal = 16'b0000001001000011;
            15'd3774: log10_cal = 16'b0000001001000100;
            15'd3775: log10_cal = 16'b0000001001000100;
            15'd3776: log10_cal = 16'b0000001001000100;
            15'd3777: log10_cal = 16'b0000001001000100;
            15'd3778: log10_cal = 16'b0000001001000100;
            15'd3779: log10_cal = 16'b0000001001000100;
            15'd3780: log10_cal = 16'b0000001001000100;
            15'd3781: log10_cal = 16'b0000001001000100;
            15'd3782: log10_cal = 16'b0000001001000101;
            15'd3783: log10_cal = 16'b0000001001000101;
            15'd3784: log10_cal = 16'b0000001001000101;
            15'd3785: log10_cal = 16'b0000001001000101;
            15'd3786: log10_cal = 16'b0000001001000101;
            15'd3787: log10_cal = 16'b0000001001000101;
            15'd3788: log10_cal = 16'b0000001001000101;
            15'd3789: log10_cal = 16'b0000001001000101;
            15'd3790: log10_cal = 16'b0000001001000101;
            15'd3791: log10_cal = 16'b0000001001000110;
            15'd3792: log10_cal = 16'b0000001001000110;
            15'd3793: log10_cal = 16'b0000001001000110;
            15'd3794: log10_cal = 16'b0000001001000110;
            15'd3795: log10_cal = 16'b0000001001000110;
            15'd3796: log10_cal = 16'b0000001001000110;
            15'd3797: log10_cal = 16'b0000001001000110;
            15'd3798: log10_cal = 16'b0000001001000110;
            15'd3799: log10_cal = 16'b0000001001000111;
            15'd3800: log10_cal = 16'b0000001001000111;
            15'd3801: log10_cal = 16'b0000001001000111;
            15'd3802: log10_cal = 16'b0000001001000111;
            15'd3803: log10_cal = 16'b0000001001000111;
            15'd3804: log10_cal = 16'b0000001001000111;
            15'd3805: log10_cal = 16'b0000001001000111;
            15'd3806: log10_cal = 16'b0000001001000111;
            15'd3807: log10_cal = 16'b0000001001000111;
            15'd3808: log10_cal = 16'b0000001001001000;
            15'd3809: log10_cal = 16'b0000001001001000;
            15'd3810: log10_cal = 16'b0000001001001000;
            15'd3811: log10_cal = 16'b0000001001001000;
            15'd3812: log10_cal = 16'b0000001001001000;
            15'd3813: log10_cal = 16'b0000001001001000;
            15'd3814: log10_cal = 16'b0000001001001000;
            15'd3815: log10_cal = 16'b0000001001001000;
            15'd3816: log10_cal = 16'b0000001001001001;
            15'd3817: log10_cal = 16'b0000001001001001;
            15'd3818: log10_cal = 16'b0000001001001001;
            15'd3819: log10_cal = 16'b0000001001001001;
            15'd3820: log10_cal = 16'b0000001001001001;
            15'd3821: log10_cal = 16'b0000001001001001;
            15'd3822: log10_cal = 16'b0000001001001001;
            15'd3823: log10_cal = 16'b0000001001001001;
            15'd3824: log10_cal = 16'b0000001001001001;
            15'd3825: log10_cal = 16'b0000001001001010;
            15'd3826: log10_cal = 16'b0000001001001010;
            15'd3827: log10_cal = 16'b0000001001001010;
            15'd3828: log10_cal = 16'b0000001001001010;
            15'd3829: log10_cal = 16'b0000001001001010;
            15'd3830: log10_cal = 16'b0000001001001010;
            15'd3831: log10_cal = 16'b0000001001001010;
            15'd3832: log10_cal = 16'b0000001001001010;
            15'd3833: log10_cal = 16'b0000001001001010;
            15'd3834: log10_cal = 16'b0000001001001011;
            15'd3835: log10_cal = 16'b0000001001001011;
            15'd3836: log10_cal = 16'b0000001001001011;
            15'd3837: log10_cal = 16'b0000001001001011;
            15'd3838: log10_cal = 16'b0000001001001011;
            15'd3839: log10_cal = 16'b0000001001001011;
            15'd3840: log10_cal = 16'b0000001001001011;
            15'd3841: log10_cal = 16'b0000001001001011;
            15'd3842: log10_cal = 16'b0000001001001100;
            15'd3843: log10_cal = 16'b0000001001001100;
            15'd3844: log10_cal = 16'b0000001001001100;
            15'd3845: log10_cal = 16'b0000001001001100;
            15'd3846: log10_cal = 16'b0000001001001100;
            15'd3847: log10_cal = 16'b0000001001001100;
            15'd3848: log10_cal = 16'b0000001001001100;
            15'd3849: log10_cal = 16'b0000001001001100;
            15'd3850: log10_cal = 16'b0000001001001100;
            15'd3851: log10_cal = 16'b0000001001001101;
            15'd3852: log10_cal = 16'b0000001001001101;
            15'd3853: log10_cal = 16'b0000001001001101;
            15'd3854: log10_cal = 16'b0000001001001101;
            15'd3855: log10_cal = 16'b0000001001001101;
            15'd3856: log10_cal = 16'b0000001001001101;
            15'd3857: log10_cal = 16'b0000001001001101;
            15'd3858: log10_cal = 16'b0000001001001101;
            15'd3859: log10_cal = 16'b0000001001001110;
            15'd3860: log10_cal = 16'b0000001001001110;
            15'd3861: log10_cal = 16'b0000001001001110;
            15'd3862: log10_cal = 16'b0000001001001110;
            15'd3863: log10_cal = 16'b0000001001001110;
            15'd3864: log10_cal = 16'b0000001001001110;
            15'd3865: log10_cal = 16'b0000001001001110;
            15'd3866: log10_cal = 16'b0000001001001110;
            15'd3867: log10_cal = 16'b0000001001001110;
            15'd3868: log10_cal = 16'b0000001001001111;
            15'd3869: log10_cal = 16'b0000001001001111;
            15'd3870: log10_cal = 16'b0000001001001111;
            15'd3871: log10_cal = 16'b0000001001001111;
            15'd3872: log10_cal = 16'b0000001001001111;
            15'd3873: log10_cal = 16'b0000001001001111;
            15'd3874: log10_cal = 16'b0000001001001111;
            15'd3875: log10_cal = 16'b0000001001001111;
            15'd3876: log10_cal = 16'b0000001001001111;
            15'd3877: log10_cal = 16'b0000001001010000;
            15'd3878: log10_cal = 16'b0000001001010000;
            15'd3879: log10_cal = 16'b0000001001010000;
            15'd3880: log10_cal = 16'b0000001001010000;
            15'd3881: log10_cal = 16'b0000001001010000;
            15'd3882: log10_cal = 16'b0000001001010000;
            15'd3883: log10_cal = 16'b0000001001010000;
            15'd3884: log10_cal = 16'b0000001001010000;
            15'd3885: log10_cal = 16'b0000001001010000;
            15'd3886: log10_cal = 16'b0000001001010001;
            15'd3887: log10_cal = 16'b0000001001010001;
            15'd3888: log10_cal = 16'b0000001001010001;
            15'd3889: log10_cal = 16'b0000001001010001;
            15'd3890: log10_cal = 16'b0000001001010001;
            15'd3891: log10_cal = 16'b0000001001010001;
            15'd3892: log10_cal = 16'b0000001001010001;
            15'd3893: log10_cal = 16'b0000001001010001;
            15'd3894: log10_cal = 16'b0000001001010010;
            15'd3895: log10_cal = 16'b0000001001010010;
            15'd3896: log10_cal = 16'b0000001001010010;
            15'd3897: log10_cal = 16'b0000001001010010;
            15'd3898: log10_cal = 16'b0000001001010010;
            15'd3899: log10_cal = 16'b0000001001010010;
            15'd3900: log10_cal = 16'b0000001001010010;
            15'd3901: log10_cal = 16'b0000001001010010;
            15'd3902: log10_cal = 16'b0000001001010010;
            15'd3903: log10_cal = 16'b0000001001010011;
            15'd3904: log10_cal = 16'b0000001001010011;
            15'd3905: log10_cal = 16'b0000001001010011;
            15'd3906: log10_cal = 16'b0000001001010011;
            15'd3907: log10_cal = 16'b0000001001010011;
            15'd3908: log10_cal = 16'b0000001001010011;
            15'd3909: log10_cal = 16'b0000001001010011;
            15'd3910: log10_cal = 16'b0000001001010011;
            15'd3911: log10_cal = 16'b0000001001010011;
            15'd3912: log10_cal = 16'b0000001001010100;
            15'd3913: log10_cal = 16'b0000001001010100;
            15'd3914: log10_cal = 16'b0000001001010100;
            15'd3915: log10_cal = 16'b0000001001010100;
            15'd3916: log10_cal = 16'b0000001001010100;
            15'd3917: log10_cal = 16'b0000001001010100;
            15'd3918: log10_cal = 16'b0000001001010100;
            15'd3919: log10_cal = 16'b0000001001010100;
            15'd3920: log10_cal = 16'b0000001001010100;
            15'd3921: log10_cal = 16'b0000001001010101;
            15'd3922: log10_cal = 16'b0000001001010101;
            15'd3923: log10_cal = 16'b0000001001010101;
            15'd3924: log10_cal = 16'b0000001001010101;
            15'd3925: log10_cal = 16'b0000001001010101;
            15'd3926: log10_cal = 16'b0000001001010101;
            15'd3927: log10_cal = 16'b0000001001010101;
            15'd3928: log10_cal = 16'b0000001001010101;
            15'd3929: log10_cal = 16'b0000001001010101;
            15'd3930: log10_cal = 16'b0000001001010110;
            15'd3931: log10_cal = 16'b0000001001010110;
            15'd3932: log10_cal = 16'b0000001001010110;
            15'd3933: log10_cal = 16'b0000001001010110;
            15'd3934: log10_cal = 16'b0000001001010110;
            15'd3935: log10_cal = 16'b0000001001010110;
            15'd3936: log10_cal = 16'b0000001001010110;
            15'd3937: log10_cal = 16'b0000001001010110;
            15'd3938: log10_cal = 16'b0000001001010111;
            15'd3939: log10_cal = 16'b0000001001010111;
            15'd3940: log10_cal = 16'b0000001001010111;
            15'd3941: log10_cal = 16'b0000001001010111;
            15'd3942: log10_cal = 16'b0000001001010111;
            15'd3943: log10_cal = 16'b0000001001010111;
            15'd3944: log10_cal = 16'b0000001001010111;
            15'd3945: log10_cal = 16'b0000001001010111;
            15'd3946: log10_cal = 16'b0000001001010111;
            15'd3947: log10_cal = 16'b0000001001011000;
            15'd3948: log10_cal = 16'b0000001001011000;
            15'd3949: log10_cal = 16'b0000001001011000;
            15'd3950: log10_cal = 16'b0000001001011000;
            15'd3951: log10_cal = 16'b0000001001011000;
            15'd3952: log10_cal = 16'b0000001001011000;
            15'd3953: log10_cal = 16'b0000001001011000;
            15'd3954: log10_cal = 16'b0000001001011000;
            15'd3955: log10_cal = 16'b0000001001011000;
            15'd3956: log10_cal = 16'b0000001001011001;
            15'd3957: log10_cal = 16'b0000001001011001;
            15'd3958: log10_cal = 16'b0000001001011001;
            15'd3959: log10_cal = 16'b0000001001011001;
            15'd3960: log10_cal = 16'b0000001001011001;
            15'd3961: log10_cal = 16'b0000001001011001;
            15'd3962: log10_cal = 16'b0000001001011001;
            15'd3963: log10_cal = 16'b0000001001011001;
            15'd3964: log10_cal = 16'b0000001001011001;
            15'd3965: log10_cal = 16'b0000001001011010;
            15'd3966: log10_cal = 16'b0000001001011010;
            15'd3967: log10_cal = 16'b0000001001011010;
            15'd3968: log10_cal = 16'b0000001001011010;
            15'd3969: log10_cal = 16'b0000001001011010;
            15'd3970: log10_cal = 16'b0000001001011010;
            15'd3971: log10_cal = 16'b0000001001011010;
            15'd3972: log10_cal = 16'b0000001001011010;
            15'd3973: log10_cal = 16'b0000001001011010;
            15'd3974: log10_cal = 16'b0000001001011011;
            15'd3975: log10_cal = 16'b0000001001011011;
            15'd3976: log10_cal = 16'b0000001001011011;
            15'd3977: log10_cal = 16'b0000001001011011;
            15'd3978: log10_cal = 16'b0000001001011011;
            15'd3979: log10_cal = 16'b0000001001011011;
            15'd3980: log10_cal = 16'b0000001001011011;
            15'd3981: log10_cal = 16'b0000001001011011;
            15'd3982: log10_cal = 16'b0000001001011011;
            15'd3983: log10_cal = 16'b0000001001011100;
            15'd3984: log10_cal = 16'b0000001001011100;
            15'd3985: log10_cal = 16'b0000001001011100;
            15'd3986: log10_cal = 16'b0000001001011100;
            15'd3987: log10_cal = 16'b0000001001011100;
            15'd3988: log10_cal = 16'b0000001001011100;
            15'd3989: log10_cal = 16'b0000001001011100;
            15'd3990: log10_cal = 16'b0000001001011100;
            15'd3991: log10_cal = 16'b0000001001011100;
            15'd3992: log10_cal = 16'b0000001001011101;
            15'd3993: log10_cal = 16'b0000001001011101;
            15'd3994: log10_cal = 16'b0000001001011101;
            15'd3995: log10_cal = 16'b0000001001011101;
            15'd3996: log10_cal = 16'b0000001001011101;
            15'd3997: log10_cal = 16'b0000001001011101;
            15'd3998: log10_cal = 16'b0000001001011101;
            15'd3999: log10_cal = 16'b0000001001011101;
            15'd4000: log10_cal = 16'b0000001001011101;
            15'd4001: log10_cal = 16'b0000001001011110;
            15'd4002: log10_cal = 16'b0000001001011110;
            15'd4003: log10_cal = 16'b0000001001011110;
            15'd4004: log10_cal = 16'b0000001001011110;
            15'd4005: log10_cal = 16'b0000001001011110;
            15'd4006: log10_cal = 16'b0000001001011110;
            15'd4007: log10_cal = 16'b0000001001011110;
            15'd4008: log10_cal = 16'b0000001001011110;
            15'd4009: log10_cal = 16'b0000001001011110;
            15'd4010: log10_cal = 16'b0000001001011111;
            15'd4011: log10_cal = 16'b0000001001011111;
            15'd4012: log10_cal = 16'b0000001001011111;
            15'd4013: log10_cal = 16'b0000001001011111;
            15'd4014: log10_cal = 16'b0000001001011111;
            15'd4015: log10_cal = 16'b0000001001011111;
            15'd4016: log10_cal = 16'b0000001001011111;
            15'd4017: log10_cal = 16'b0000001001011111;
            15'd4018: log10_cal = 16'b0000001001011111;
            15'd4019: log10_cal = 16'b0000001001100000;
            15'd4020: log10_cal = 16'b0000001001100000;
            15'd4021: log10_cal = 16'b0000001001100000;
            15'd4022: log10_cal = 16'b0000001001100000;
            15'd4023: log10_cal = 16'b0000001001100000;
            15'd4024: log10_cal = 16'b0000001001100000;
            15'd4025: log10_cal = 16'b0000001001100000;
            15'd4026: log10_cal = 16'b0000001001100000;
            15'd4027: log10_cal = 16'b0000001001100000;
            15'd4028: log10_cal = 16'b0000001001100001;
            15'd4029: log10_cal = 16'b0000001001100001;
            15'd4030: log10_cal = 16'b0000001001100001;
            15'd4031: log10_cal = 16'b0000001001100001;
            15'd4032: log10_cal = 16'b0000001001100001;
            15'd4033: log10_cal = 16'b0000001001100001;
            15'd4034: log10_cal = 16'b0000001001100001;
            15'd4035: log10_cal = 16'b0000001001100001;
            15'd4036: log10_cal = 16'b0000001001100001;
            15'd4037: log10_cal = 16'b0000001001100010;
            15'd4038: log10_cal = 16'b0000001001100010;
            15'd4039: log10_cal = 16'b0000001001100010;
            15'd4040: log10_cal = 16'b0000001001100010;
            15'd4041: log10_cal = 16'b0000001001100010;
            15'd4042: log10_cal = 16'b0000001001100010;
            15'd4043: log10_cal = 16'b0000001001100010;
            15'd4044: log10_cal = 16'b0000001001100010;
            15'd4045: log10_cal = 16'b0000001001100010;
            15'd4046: log10_cal = 16'b0000001001100011;
            15'd4047: log10_cal = 16'b0000001001100011;
            15'd4048: log10_cal = 16'b0000001001100011;
            15'd4049: log10_cal = 16'b0000001001100011;
            15'd4050: log10_cal = 16'b0000001001100011;
            15'd4051: log10_cal = 16'b0000001001100011;
            15'd4052: log10_cal = 16'b0000001001100011;
            15'd4053: log10_cal = 16'b0000001001100011;
            15'd4054: log10_cal = 16'b0000001001100011;
            15'd4055: log10_cal = 16'b0000001001100100;
            15'd4056: log10_cal = 16'b0000001001100100;
            15'd4057: log10_cal = 16'b0000001001100100;
            15'd4058: log10_cal = 16'b0000001001100100;
            15'd4059: log10_cal = 16'b0000001001100100;
            15'd4060: log10_cal = 16'b0000001001100100;
            15'd4061: log10_cal = 16'b0000001001100100;
            15'd4062: log10_cal = 16'b0000001001100100;
            15'd4063: log10_cal = 16'b0000001001100100;
            15'd4064: log10_cal = 16'b0000001001100101;
            15'd4065: log10_cal = 16'b0000001001100101;
            15'd4066: log10_cal = 16'b0000001001100101;
            15'd4067: log10_cal = 16'b0000001001100101;
            15'd4068: log10_cal = 16'b0000001001100101;
            15'd4069: log10_cal = 16'b0000001001100101;
            15'd4070: log10_cal = 16'b0000001001100101;
            15'd4071: log10_cal = 16'b0000001001100101;
            15'd4072: log10_cal = 16'b0000001001100101;
            15'd4073: log10_cal = 16'b0000001001100110;
            15'd4074: log10_cal = 16'b0000001001100110;
            15'd4075: log10_cal = 16'b0000001001100110;
            15'd4076: log10_cal = 16'b0000001001100110;
            15'd4077: log10_cal = 16'b0000001001100110;
            15'd4078: log10_cal = 16'b0000001001100110;
            15'd4079: log10_cal = 16'b0000001001100110;
            15'd4080: log10_cal = 16'b0000001001100110;
            15'd4081: log10_cal = 16'b0000001001100110;
            15'd4082: log10_cal = 16'b0000001001100110;
            15'd4083: log10_cal = 16'b0000001001100111;
            15'd4084: log10_cal = 16'b0000001001100111;
            15'd4085: log10_cal = 16'b0000001001100111;
            15'd4086: log10_cal = 16'b0000001001100111;
            15'd4087: log10_cal = 16'b0000001001100111;
            15'd4088: log10_cal = 16'b0000001001100111;
            15'd4089: log10_cal = 16'b0000001001100111;
            15'd4090: log10_cal = 16'b0000001001100111;
            15'd4091: log10_cal = 16'b0000001001100111;
            15'd4092: log10_cal = 16'b0000001001101000;
            15'd4093: log10_cal = 16'b0000001001101000;
            15'd4094: log10_cal = 16'b0000001001101000;
            15'd4095: log10_cal = 16'b0000001001101000;
            15'd4096: log10_cal = 16'b0000001001101000;
            15'd4097: log10_cal = 16'b0000001001101000;
            15'd4098: log10_cal = 16'b0000001001101000;
            15'd4099: log10_cal = 16'b0000001001101000;
            15'd4100: log10_cal = 16'b0000001001101000;
            15'd4101: log10_cal = 16'b0000001001101001;
            15'd4102: log10_cal = 16'b0000001001101001;
            15'd4103: log10_cal = 16'b0000001001101001;
            15'd4104: log10_cal = 16'b0000001001101001;
            15'd4105: log10_cal = 16'b0000001001101001;
            15'd4106: log10_cal = 16'b0000001001101001;
            15'd4107: log10_cal = 16'b0000001001101001;
            15'd4108: log10_cal = 16'b0000001001101001;
            15'd4109: log10_cal = 16'b0000001001101001;
            15'd4110: log10_cal = 16'b0000001001101010;
            15'd4111: log10_cal = 16'b0000001001101010;
            15'd4112: log10_cal = 16'b0000001001101010;
            15'd4113: log10_cal = 16'b0000001001101010;
            15'd4114: log10_cal = 16'b0000001001101010;
            15'd4115: log10_cal = 16'b0000001001101010;
            15'd4116: log10_cal = 16'b0000001001101010;
            15'd4117: log10_cal = 16'b0000001001101010;
            15'd4118: log10_cal = 16'b0000001001101010;
            15'd4119: log10_cal = 16'b0000001001101010;
            15'd4120: log10_cal = 16'b0000001001101011;
            15'd4121: log10_cal = 16'b0000001001101011;
            15'd4122: log10_cal = 16'b0000001001101011;
            15'd4123: log10_cal = 16'b0000001001101011;
            15'd4124: log10_cal = 16'b0000001001101011;
            15'd4125: log10_cal = 16'b0000001001101011;
            15'd4126: log10_cal = 16'b0000001001101011;
            15'd4127: log10_cal = 16'b0000001001101011;
            15'd4128: log10_cal = 16'b0000001001101011;
            15'd4129: log10_cal = 16'b0000001001101100;
            15'd4130: log10_cal = 16'b0000001001101100;
            15'd4131: log10_cal = 16'b0000001001101100;
            15'd4132: log10_cal = 16'b0000001001101100;
            15'd4133: log10_cal = 16'b0000001001101100;
            15'd4134: log10_cal = 16'b0000001001101100;
            15'd4135: log10_cal = 16'b0000001001101100;
            15'd4136: log10_cal = 16'b0000001001101100;
            15'd4137: log10_cal = 16'b0000001001101100;
            15'd4138: log10_cal = 16'b0000001001101101;
            15'd4139: log10_cal = 16'b0000001001101101;
            15'd4140: log10_cal = 16'b0000001001101101;
            15'd4141: log10_cal = 16'b0000001001101101;
            15'd4142: log10_cal = 16'b0000001001101101;
            15'd4143: log10_cal = 16'b0000001001101101;
            15'd4144: log10_cal = 16'b0000001001101101;
            15'd4145: log10_cal = 16'b0000001001101101;
            15'd4146: log10_cal = 16'b0000001001101101;
            15'd4147: log10_cal = 16'b0000001001101110;
            15'd4148: log10_cal = 16'b0000001001101110;
            15'd4149: log10_cal = 16'b0000001001101110;
            15'd4150: log10_cal = 16'b0000001001101110;
            15'd4151: log10_cal = 16'b0000001001101110;
            15'd4152: log10_cal = 16'b0000001001101110;
            15'd4153: log10_cal = 16'b0000001001101110;
            15'd4154: log10_cal = 16'b0000001001101110;
            15'd4155: log10_cal = 16'b0000001001101110;
            15'd4156: log10_cal = 16'b0000001001101110;
            15'd4157: log10_cal = 16'b0000001001101111;
            15'd4158: log10_cal = 16'b0000001001101111;
            15'd4159: log10_cal = 16'b0000001001101111;
            15'd4160: log10_cal = 16'b0000001001101111;
            15'd4161: log10_cal = 16'b0000001001101111;
            15'd4162: log10_cal = 16'b0000001001101111;
            15'd4163: log10_cal = 16'b0000001001101111;
            15'd4164: log10_cal = 16'b0000001001101111;
            15'd4165: log10_cal = 16'b0000001001101111;
            15'd4166: log10_cal = 16'b0000001001110000;
            15'd4167: log10_cal = 16'b0000001001110000;
            15'd4168: log10_cal = 16'b0000001001110000;
            15'd4169: log10_cal = 16'b0000001001110000;
            15'd4170: log10_cal = 16'b0000001001110000;
            15'd4171: log10_cal = 16'b0000001001110000;
            15'd4172: log10_cal = 16'b0000001001110000;
            15'd4173: log10_cal = 16'b0000001001110000;
            15'd4174: log10_cal = 16'b0000001001110000;
            15'd4175: log10_cal = 16'b0000001001110001;
            15'd4176: log10_cal = 16'b0000001001110001;
            15'd4177: log10_cal = 16'b0000001001110001;
            15'd4178: log10_cal = 16'b0000001001110001;
            15'd4179: log10_cal = 16'b0000001001110001;
            15'd4180: log10_cal = 16'b0000001001110001;
            15'd4181: log10_cal = 16'b0000001001110001;
            15'd4182: log10_cal = 16'b0000001001110001;
            15'd4183: log10_cal = 16'b0000001001110001;
            15'd4184: log10_cal = 16'b0000001001110001;
            15'd4185: log10_cal = 16'b0000001001110010;
            15'd4186: log10_cal = 16'b0000001001110010;
            15'd4187: log10_cal = 16'b0000001001110010;
            15'd4188: log10_cal = 16'b0000001001110010;
            15'd4189: log10_cal = 16'b0000001001110010;
            15'd4190: log10_cal = 16'b0000001001110010;
            15'd4191: log10_cal = 16'b0000001001110010;
            15'd4192: log10_cal = 16'b0000001001110010;
            15'd4193: log10_cal = 16'b0000001001110010;
            15'd4194: log10_cal = 16'b0000001001110011;
            15'd4195: log10_cal = 16'b0000001001110011;
            15'd4196: log10_cal = 16'b0000001001110011;
            15'd4197: log10_cal = 16'b0000001001110011;
            15'd4198: log10_cal = 16'b0000001001110011;
            15'd4199: log10_cal = 16'b0000001001110011;
            15'd4200: log10_cal = 16'b0000001001110011;
            15'd4201: log10_cal = 16'b0000001001110011;
            15'd4202: log10_cal = 16'b0000001001110011;
            15'd4203: log10_cal = 16'b0000001001110011;
            15'd4204: log10_cal = 16'b0000001001110100;
            15'd4205: log10_cal = 16'b0000001001110100;
            15'd4206: log10_cal = 16'b0000001001110100;
            15'd4207: log10_cal = 16'b0000001001110100;
            15'd4208: log10_cal = 16'b0000001001110100;
            15'd4209: log10_cal = 16'b0000001001110100;
            15'd4210: log10_cal = 16'b0000001001110100;
            15'd4211: log10_cal = 16'b0000001001110100;
            15'd4212: log10_cal = 16'b0000001001110100;
            15'd4213: log10_cal = 16'b0000001001110101;
            15'd4214: log10_cal = 16'b0000001001110101;
            15'd4215: log10_cal = 16'b0000001001110101;
            15'd4216: log10_cal = 16'b0000001001110101;
            15'd4217: log10_cal = 16'b0000001001110101;
            15'd4218: log10_cal = 16'b0000001001110101;
            15'd4219: log10_cal = 16'b0000001001110101;
            15'd4220: log10_cal = 16'b0000001001110101;
            15'd4221: log10_cal = 16'b0000001001110101;
            15'd4222: log10_cal = 16'b0000001001110101;
            15'd4223: log10_cal = 16'b0000001001110110;
            15'd4224: log10_cal = 16'b0000001001110110;
            15'd4225: log10_cal = 16'b0000001001110110;
            15'd4226: log10_cal = 16'b0000001001110110;
            15'd4227: log10_cal = 16'b0000001001110110;
            15'd4228: log10_cal = 16'b0000001001110110;
            15'd4229: log10_cal = 16'b0000001001110110;
            15'd4230: log10_cal = 16'b0000001001110110;
            15'd4231: log10_cal = 16'b0000001001110110;
            15'd4232: log10_cal = 16'b0000001001110111;
            15'd4233: log10_cal = 16'b0000001001110111;
            15'd4234: log10_cal = 16'b0000001001110111;
            15'd4235: log10_cal = 16'b0000001001110111;
            15'd4236: log10_cal = 16'b0000001001110111;
            15'd4237: log10_cal = 16'b0000001001110111;
            15'd4238: log10_cal = 16'b0000001001110111;
            15'd4239: log10_cal = 16'b0000001001110111;
            15'd4240: log10_cal = 16'b0000001001110111;
            15'd4241: log10_cal = 16'b0000001001110111;
            15'd4242: log10_cal = 16'b0000001001111000;
            15'd4243: log10_cal = 16'b0000001001111000;
            15'd4244: log10_cal = 16'b0000001001111000;
            15'd4245: log10_cal = 16'b0000001001111000;
            15'd4246: log10_cal = 16'b0000001001111000;
            15'd4247: log10_cal = 16'b0000001001111000;
            15'd4248: log10_cal = 16'b0000001001111000;
            15'd4249: log10_cal = 16'b0000001001111000;
            15'd4250: log10_cal = 16'b0000001001111000;
            15'd4251: log10_cal = 16'b0000001001111001;
            15'd4252: log10_cal = 16'b0000001001111001;
            15'd4253: log10_cal = 16'b0000001001111001;
            15'd4254: log10_cal = 16'b0000001001111001;
            15'd4255: log10_cal = 16'b0000001001111001;
            15'd4256: log10_cal = 16'b0000001001111001;
            15'd4257: log10_cal = 16'b0000001001111001;
            15'd4258: log10_cal = 16'b0000001001111001;
            15'd4259: log10_cal = 16'b0000001001111001;
            15'd4260: log10_cal = 16'b0000001001111001;
            15'd4261: log10_cal = 16'b0000001001111010;
            15'd4262: log10_cal = 16'b0000001001111010;
            15'd4263: log10_cal = 16'b0000001001111010;
            15'd4264: log10_cal = 16'b0000001001111010;
            15'd4265: log10_cal = 16'b0000001001111010;
            15'd4266: log10_cal = 16'b0000001001111010;
            15'd4267: log10_cal = 16'b0000001001111010;
            15'd4268: log10_cal = 16'b0000001001111010;
            15'd4269: log10_cal = 16'b0000001001111010;
            15'd4270: log10_cal = 16'b0000001001111011;
            15'd4271: log10_cal = 16'b0000001001111011;
            15'd4272: log10_cal = 16'b0000001001111011;
            15'd4273: log10_cal = 16'b0000001001111011;
            15'd4274: log10_cal = 16'b0000001001111011;
            15'd4275: log10_cal = 16'b0000001001111011;
            15'd4276: log10_cal = 16'b0000001001111011;
            15'd4277: log10_cal = 16'b0000001001111011;
            15'd4278: log10_cal = 16'b0000001001111011;
            15'd4279: log10_cal = 16'b0000001001111011;
            15'd4280: log10_cal = 16'b0000001001111100;
            15'd4281: log10_cal = 16'b0000001001111100;
            15'd4282: log10_cal = 16'b0000001001111100;
            15'd4283: log10_cal = 16'b0000001001111100;
            15'd4284: log10_cal = 16'b0000001001111100;
            15'd4285: log10_cal = 16'b0000001001111100;
            15'd4286: log10_cal = 16'b0000001001111100;
            15'd4287: log10_cal = 16'b0000001001111100;
            15'd4288: log10_cal = 16'b0000001001111100;
            15'd4289: log10_cal = 16'b0000001001111100;
            15'd4290: log10_cal = 16'b0000001001111101;
            15'd4291: log10_cal = 16'b0000001001111101;
            15'd4292: log10_cal = 16'b0000001001111101;
            15'd4293: log10_cal = 16'b0000001001111101;
            15'd4294: log10_cal = 16'b0000001001111101;
            15'd4295: log10_cal = 16'b0000001001111101;
            15'd4296: log10_cal = 16'b0000001001111101;
            15'd4297: log10_cal = 16'b0000001001111101;
            15'd4298: log10_cal = 16'b0000001001111101;
            15'd4299: log10_cal = 16'b0000001001111110;
            15'd4300: log10_cal = 16'b0000001001111110;
            15'd4301: log10_cal = 16'b0000001001111110;
            15'd4302: log10_cal = 16'b0000001001111110;
            15'd4303: log10_cal = 16'b0000001001111110;
            15'd4304: log10_cal = 16'b0000001001111110;
            15'd4305: log10_cal = 16'b0000001001111110;
            15'd4306: log10_cal = 16'b0000001001111110;
            15'd4307: log10_cal = 16'b0000001001111110;
            15'd4308: log10_cal = 16'b0000001001111110;
            15'd4309: log10_cal = 16'b0000001001111111;
            15'd4310: log10_cal = 16'b0000001001111111;
            15'd4311: log10_cal = 16'b0000001001111111;
            15'd4312: log10_cal = 16'b0000001001111111;
            15'd4313: log10_cal = 16'b0000001001111111;
            15'd4314: log10_cal = 16'b0000001001111111;
            15'd4315: log10_cal = 16'b0000001001111111;
            15'd4316: log10_cal = 16'b0000001001111111;
            15'd4317: log10_cal = 16'b0000001001111111;
            15'd4318: log10_cal = 16'b0000001001111111;
            15'd4319: log10_cal = 16'b0000001010000000;
            15'd4320: log10_cal = 16'b0000001010000000;
            15'd4321: log10_cal = 16'b0000001010000000;
            15'd4322: log10_cal = 16'b0000001010000000;
            15'd4323: log10_cal = 16'b0000001010000000;
            15'd4324: log10_cal = 16'b0000001010000000;
            15'd4325: log10_cal = 16'b0000001010000000;
            15'd4326: log10_cal = 16'b0000001010000000;
            15'd4327: log10_cal = 16'b0000001010000000;
            15'd4328: log10_cal = 16'b0000001010000001;
            15'd4329: log10_cal = 16'b0000001010000001;
            15'd4330: log10_cal = 16'b0000001010000001;
            15'd4331: log10_cal = 16'b0000001010000001;
            15'd4332: log10_cal = 16'b0000001010000001;
            15'd4333: log10_cal = 16'b0000001010000001;
            15'd4334: log10_cal = 16'b0000001010000001;
            15'd4335: log10_cal = 16'b0000001010000001;
            15'd4336: log10_cal = 16'b0000001010000001;
            15'd4337: log10_cal = 16'b0000001010000001;
            15'd4338: log10_cal = 16'b0000001010000010;
            15'd4339: log10_cal = 16'b0000001010000010;
            15'd4340: log10_cal = 16'b0000001010000010;
            15'd4341: log10_cal = 16'b0000001010000010;
            15'd4342: log10_cal = 16'b0000001010000010;
            15'd4343: log10_cal = 16'b0000001010000010;
            15'd4344: log10_cal = 16'b0000001010000010;
            15'd4345: log10_cal = 16'b0000001010000010;
            15'd4346: log10_cal = 16'b0000001010000010;
            15'd4347: log10_cal = 16'b0000001010000010;
            15'd4348: log10_cal = 16'b0000001010000011;
            15'd4349: log10_cal = 16'b0000001010000011;
            15'd4350: log10_cal = 16'b0000001010000011;
            15'd4351: log10_cal = 16'b0000001010000011;
            15'd4352: log10_cal = 16'b0000001010000011;
            15'd4353: log10_cal = 16'b0000001010000011;
            15'd4354: log10_cal = 16'b0000001010000011;
            15'd4355: log10_cal = 16'b0000001010000011;
            15'd4356: log10_cal = 16'b0000001010000011;
            15'd4357: log10_cal = 16'b0000001010000011;
            15'd4358: log10_cal = 16'b0000001010000100;
            15'd4359: log10_cal = 16'b0000001010000100;
            15'd4360: log10_cal = 16'b0000001010000100;
            15'd4361: log10_cal = 16'b0000001010000100;
            15'd4362: log10_cal = 16'b0000001010000100;
            15'd4363: log10_cal = 16'b0000001010000100;
            15'd4364: log10_cal = 16'b0000001010000100;
            15'd4365: log10_cal = 16'b0000001010000100;
            15'd4366: log10_cal = 16'b0000001010000100;
            15'd4367: log10_cal = 16'b0000001010000101;
            15'd4368: log10_cal = 16'b0000001010000101;
            15'd4369: log10_cal = 16'b0000001010000101;
            15'd4370: log10_cal = 16'b0000001010000101;
            15'd4371: log10_cal = 16'b0000001010000101;
            15'd4372: log10_cal = 16'b0000001010000101;
            15'd4373: log10_cal = 16'b0000001010000101;
            15'd4374: log10_cal = 16'b0000001010000101;
            15'd4375: log10_cal = 16'b0000001010000101;
            15'd4376: log10_cal = 16'b0000001010000101;
            15'd4377: log10_cal = 16'b0000001010000110;
            15'd4378: log10_cal = 16'b0000001010000110;
            15'd4379: log10_cal = 16'b0000001010000110;
            15'd4380: log10_cal = 16'b0000001010000110;
            15'd4381: log10_cal = 16'b0000001010000110;
            15'd4382: log10_cal = 16'b0000001010000110;
            15'd4383: log10_cal = 16'b0000001010000110;
            15'd4384: log10_cal = 16'b0000001010000110;
            15'd4385: log10_cal = 16'b0000001010000110;
            15'd4386: log10_cal = 16'b0000001010000110;
            15'd4387: log10_cal = 16'b0000001010000111;
            15'd4388: log10_cal = 16'b0000001010000111;
            15'd4389: log10_cal = 16'b0000001010000111;
            15'd4390: log10_cal = 16'b0000001010000111;
            15'd4391: log10_cal = 16'b0000001010000111;
            15'd4392: log10_cal = 16'b0000001010000111;
            15'd4393: log10_cal = 16'b0000001010000111;
            15'd4394: log10_cal = 16'b0000001010000111;
            15'd4395: log10_cal = 16'b0000001010000111;
            15'd4396: log10_cal = 16'b0000001010000111;
            15'd4397: log10_cal = 16'b0000001010001000;
            15'd4398: log10_cal = 16'b0000001010001000;
            15'd4399: log10_cal = 16'b0000001010001000;
            15'd4400: log10_cal = 16'b0000001010001000;
            15'd4401: log10_cal = 16'b0000001010001000;
            15'd4402: log10_cal = 16'b0000001010001000;
            15'd4403: log10_cal = 16'b0000001010001000;
            15'd4404: log10_cal = 16'b0000001010001000;
            15'd4405: log10_cal = 16'b0000001010001000;
            15'd4406: log10_cal = 16'b0000001010001000;
            15'd4407: log10_cal = 16'b0000001010001001;
            15'd4408: log10_cal = 16'b0000001010001001;
            15'd4409: log10_cal = 16'b0000001010001001;
            15'd4410: log10_cal = 16'b0000001010001001;
            15'd4411: log10_cal = 16'b0000001010001001;
            15'd4412: log10_cal = 16'b0000001010001001;
            15'd4413: log10_cal = 16'b0000001010001001;
            15'd4414: log10_cal = 16'b0000001010001001;
            15'd4415: log10_cal = 16'b0000001010001001;
            15'd4416: log10_cal = 16'b0000001010001001;
            15'd4417: log10_cal = 16'b0000001010001010;
            15'd4418: log10_cal = 16'b0000001010001010;
            15'd4419: log10_cal = 16'b0000001010001010;
            15'd4420: log10_cal = 16'b0000001010001010;
            15'd4421: log10_cal = 16'b0000001010001010;
            15'd4422: log10_cal = 16'b0000001010001010;
            15'd4423: log10_cal = 16'b0000001010001010;
            15'd4424: log10_cal = 16'b0000001010001010;
            15'd4425: log10_cal = 16'b0000001010001010;
            15'd4426: log10_cal = 16'b0000001010001010;
            15'd4427: log10_cal = 16'b0000001010001011;
            15'd4428: log10_cal = 16'b0000001010001011;
            15'd4429: log10_cal = 16'b0000001010001011;
            15'd4430: log10_cal = 16'b0000001010001011;
            15'd4431: log10_cal = 16'b0000001010001011;
            15'd4432: log10_cal = 16'b0000001010001011;
            15'd4433: log10_cal = 16'b0000001010001011;
            15'd4434: log10_cal = 16'b0000001010001011;
            15'd4435: log10_cal = 16'b0000001010001011;
            15'd4436: log10_cal = 16'b0000001010001011;
            15'd4437: log10_cal = 16'b0000001010001100;
            15'd4438: log10_cal = 16'b0000001010001100;
            15'd4439: log10_cal = 16'b0000001010001100;
            15'd4440: log10_cal = 16'b0000001010001100;
            15'd4441: log10_cal = 16'b0000001010001100;
            15'd4442: log10_cal = 16'b0000001010001100;
            15'd4443: log10_cal = 16'b0000001010001100;
            15'd4444: log10_cal = 16'b0000001010001100;
            15'd4445: log10_cal = 16'b0000001010001100;
            15'd4446: log10_cal = 16'b0000001010001100;
            15'd4447: log10_cal = 16'b0000001010001101;
            15'd4448: log10_cal = 16'b0000001010001101;
            15'd4449: log10_cal = 16'b0000001010001101;
            15'd4450: log10_cal = 16'b0000001010001101;
            15'd4451: log10_cal = 16'b0000001010001101;
            15'd4452: log10_cal = 16'b0000001010001101;
            15'd4453: log10_cal = 16'b0000001010001101;
            15'd4454: log10_cal = 16'b0000001010001101;
            15'd4455: log10_cal = 16'b0000001010001101;
            15'd4456: log10_cal = 16'b0000001010001101;
            15'd4457: log10_cal = 16'b0000001010001110;
            15'd4458: log10_cal = 16'b0000001010001110;
            15'd4459: log10_cal = 16'b0000001010001110;
            15'd4460: log10_cal = 16'b0000001010001110;
            15'd4461: log10_cal = 16'b0000001010001110;
            15'd4462: log10_cal = 16'b0000001010001110;
            15'd4463: log10_cal = 16'b0000001010001110;
            15'd4464: log10_cal = 16'b0000001010001110;
            15'd4465: log10_cal = 16'b0000001010001110;
            15'd4466: log10_cal = 16'b0000001010001110;
            15'd4467: log10_cal = 16'b0000001010001111;
            15'd4468: log10_cal = 16'b0000001010001111;
            15'd4469: log10_cal = 16'b0000001010001111;
            15'd4470: log10_cal = 16'b0000001010001111;
            15'd4471: log10_cal = 16'b0000001010001111;
            15'd4472: log10_cal = 16'b0000001010001111;
            15'd4473: log10_cal = 16'b0000001010001111;
            15'd4474: log10_cal = 16'b0000001010001111;
            15'd4475: log10_cal = 16'b0000001010001111;
            15'd4476: log10_cal = 16'b0000001010001111;
            15'd4477: log10_cal = 16'b0000001010010000;
            15'd4478: log10_cal = 16'b0000001010010000;
            15'd4479: log10_cal = 16'b0000001010010000;
            15'd4480: log10_cal = 16'b0000001010010000;
            15'd4481: log10_cal = 16'b0000001010010000;
            15'd4482: log10_cal = 16'b0000001010010000;
            15'd4483: log10_cal = 16'b0000001010010000;
            15'd4484: log10_cal = 16'b0000001010010000;
            15'd4485: log10_cal = 16'b0000001010010000;
            15'd4486: log10_cal = 16'b0000001010010000;
            15'd4487: log10_cal = 16'b0000001010010001;
            15'd4488: log10_cal = 16'b0000001010010001;
            15'd4489: log10_cal = 16'b0000001010010001;
            15'd4490: log10_cal = 16'b0000001010010001;
            15'd4491: log10_cal = 16'b0000001010010001;
            15'd4492: log10_cal = 16'b0000001010010001;
            15'd4493: log10_cal = 16'b0000001010010001;
            15'd4494: log10_cal = 16'b0000001010010001;
            15'd4495: log10_cal = 16'b0000001010010001;
            15'd4496: log10_cal = 16'b0000001010010001;
            15'd4497: log10_cal = 16'b0000001010010010;
            15'd4498: log10_cal = 16'b0000001010010010;
            15'd4499: log10_cal = 16'b0000001010010010;
            15'd4500: log10_cal = 16'b0000001010010010;
            15'd4501: log10_cal = 16'b0000001010010010;
            15'd4502: log10_cal = 16'b0000001010010010;
            15'd4503: log10_cal = 16'b0000001010010010;
            15'd4504: log10_cal = 16'b0000001010010010;
            15'd4505: log10_cal = 16'b0000001010010010;
            15'd4506: log10_cal = 16'b0000001010010010;
            15'd4507: log10_cal = 16'b0000001010010011;
            15'd4508: log10_cal = 16'b0000001010010011;
            15'd4509: log10_cal = 16'b0000001010010011;
            15'd4510: log10_cal = 16'b0000001010010011;
            15'd4511: log10_cal = 16'b0000001010010011;
            15'd4512: log10_cal = 16'b0000001010010011;
            15'd4513: log10_cal = 16'b0000001010010011;
            15'd4514: log10_cal = 16'b0000001010010011;
            15'd4515: log10_cal = 16'b0000001010010011;
            15'd4516: log10_cal = 16'b0000001010010011;
            15'd4517: log10_cal = 16'b0000001010010100;
            15'd4518: log10_cal = 16'b0000001010010100;
            15'd4519: log10_cal = 16'b0000001010010100;
            15'd4520: log10_cal = 16'b0000001010010100;
            15'd4521: log10_cal = 16'b0000001010010100;
            15'd4522: log10_cal = 16'b0000001010010100;
            15'd4523: log10_cal = 16'b0000001010010100;
            15'd4524: log10_cal = 16'b0000001010010100;
            15'd4525: log10_cal = 16'b0000001010010100;
            15'd4526: log10_cal = 16'b0000001010010100;
            15'd4527: log10_cal = 16'b0000001010010101;
            15'd4528: log10_cal = 16'b0000001010010101;
            15'd4529: log10_cal = 16'b0000001010010101;
            15'd4530: log10_cal = 16'b0000001010010101;
            15'd4531: log10_cal = 16'b0000001010010101;
            15'd4532: log10_cal = 16'b0000001010010101;
            15'd4533: log10_cal = 16'b0000001010010101;
            15'd4534: log10_cal = 16'b0000001010010101;
            15'd4535: log10_cal = 16'b0000001010010101;
            15'd4536: log10_cal = 16'b0000001010010101;
            15'd4537: log10_cal = 16'b0000001010010101;
            15'd4538: log10_cal = 16'b0000001010010110;
            15'd4539: log10_cal = 16'b0000001010010110;
            15'd4540: log10_cal = 16'b0000001010010110;
            15'd4541: log10_cal = 16'b0000001010010110;
            15'd4542: log10_cal = 16'b0000001010010110;
            15'd4543: log10_cal = 16'b0000001010010110;
            15'd4544: log10_cal = 16'b0000001010010110;
            15'd4545: log10_cal = 16'b0000001010010110;
            15'd4546: log10_cal = 16'b0000001010010110;
            15'd4547: log10_cal = 16'b0000001010010110;
            15'd4548: log10_cal = 16'b0000001010010111;
            15'd4549: log10_cal = 16'b0000001010010111;
            15'd4550: log10_cal = 16'b0000001010010111;
            15'd4551: log10_cal = 16'b0000001010010111;
            15'd4552: log10_cal = 16'b0000001010010111;
            15'd4553: log10_cal = 16'b0000001010010111;
            15'd4554: log10_cal = 16'b0000001010010111;
            15'd4555: log10_cal = 16'b0000001010010111;
            15'd4556: log10_cal = 16'b0000001010010111;
            15'd4557: log10_cal = 16'b0000001010010111;
            15'd4558: log10_cal = 16'b0000001010011000;
            15'd4559: log10_cal = 16'b0000001010011000;
            15'd4560: log10_cal = 16'b0000001010011000;
            15'd4561: log10_cal = 16'b0000001010011000;
            15'd4562: log10_cal = 16'b0000001010011000;
            15'd4563: log10_cal = 16'b0000001010011000;
            15'd4564: log10_cal = 16'b0000001010011000;
            15'd4565: log10_cal = 16'b0000001010011000;
            15'd4566: log10_cal = 16'b0000001010011000;
            15'd4567: log10_cal = 16'b0000001010011000;
            15'd4568: log10_cal = 16'b0000001010011001;
            15'd4569: log10_cal = 16'b0000001010011001;
            15'd4570: log10_cal = 16'b0000001010011001;
            15'd4571: log10_cal = 16'b0000001010011001;
            15'd4572: log10_cal = 16'b0000001010011001;
            15'd4573: log10_cal = 16'b0000001010011001;
            15'd4574: log10_cal = 16'b0000001010011001;
            15'd4575: log10_cal = 16'b0000001010011001;
            15'd4576: log10_cal = 16'b0000001010011001;
            15'd4577: log10_cal = 16'b0000001010011001;
            15'd4578: log10_cal = 16'b0000001010011001;
            15'd4579: log10_cal = 16'b0000001010011010;
            15'd4580: log10_cal = 16'b0000001010011010;
            15'd4581: log10_cal = 16'b0000001010011010;
            15'd4582: log10_cal = 16'b0000001010011010;
            15'd4583: log10_cal = 16'b0000001010011010;
            15'd4584: log10_cal = 16'b0000001010011010;
            15'd4585: log10_cal = 16'b0000001010011010;
            15'd4586: log10_cal = 16'b0000001010011010;
            15'd4587: log10_cal = 16'b0000001010011010;
            15'd4588: log10_cal = 16'b0000001010011010;
            15'd4589: log10_cal = 16'b0000001010011011;
            15'd4590: log10_cal = 16'b0000001010011011;
            15'd4591: log10_cal = 16'b0000001010011011;
            15'd4592: log10_cal = 16'b0000001010011011;
            15'd4593: log10_cal = 16'b0000001010011011;
            15'd4594: log10_cal = 16'b0000001010011011;
            15'd4595: log10_cal = 16'b0000001010011011;
            15'd4596: log10_cal = 16'b0000001010011011;
            15'd4597: log10_cal = 16'b0000001010011011;
            15'd4598: log10_cal = 16'b0000001010011011;
            15'd4599: log10_cal = 16'b0000001010011100;
            15'd4600: log10_cal = 16'b0000001010011100;
            15'd4601: log10_cal = 16'b0000001010011100;
            15'd4602: log10_cal = 16'b0000001010011100;
            15'd4603: log10_cal = 16'b0000001010011100;
            15'd4604: log10_cal = 16'b0000001010011100;
            15'd4605: log10_cal = 16'b0000001010011100;
            15'd4606: log10_cal = 16'b0000001010011100;
            15'd4607: log10_cal = 16'b0000001010011100;
            15'd4608: log10_cal = 16'b0000001010011100;
            15'd4609: log10_cal = 16'b0000001010011100;
            15'd4610: log10_cal = 16'b0000001010011101;
            15'd4611: log10_cal = 16'b0000001010011101;
            15'd4612: log10_cal = 16'b0000001010011101;
            15'd4613: log10_cal = 16'b0000001010011101;
            15'd4614: log10_cal = 16'b0000001010011101;
            15'd4615: log10_cal = 16'b0000001010011101;
            15'd4616: log10_cal = 16'b0000001010011101;
            15'd4617: log10_cal = 16'b0000001010011101;
            15'd4618: log10_cal = 16'b0000001010011101;
            15'd4619: log10_cal = 16'b0000001010011101;
            15'd4620: log10_cal = 16'b0000001010011110;
            15'd4621: log10_cal = 16'b0000001010011110;
            15'd4622: log10_cal = 16'b0000001010011110;
            15'd4623: log10_cal = 16'b0000001010011110;
            15'd4624: log10_cal = 16'b0000001010011110;
            15'd4625: log10_cal = 16'b0000001010011110;
            15'd4626: log10_cal = 16'b0000001010011110;
            15'd4627: log10_cal = 16'b0000001010011110;
            15'd4628: log10_cal = 16'b0000001010011110;
            15'd4629: log10_cal = 16'b0000001010011110;
            15'd4630: log10_cal = 16'b0000001010011111;
            15'd4631: log10_cal = 16'b0000001010011111;
            15'd4632: log10_cal = 16'b0000001010011111;
            15'd4633: log10_cal = 16'b0000001010011111;
            15'd4634: log10_cal = 16'b0000001010011111;
            15'd4635: log10_cal = 16'b0000001010011111;
            15'd4636: log10_cal = 16'b0000001010011111;
            15'd4637: log10_cal = 16'b0000001010011111;
            15'd4638: log10_cal = 16'b0000001010011111;
            15'd4639: log10_cal = 16'b0000001010011111;
            15'd4640: log10_cal = 16'b0000001010011111;
            15'd4641: log10_cal = 16'b0000001010100000;
            15'd4642: log10_cal = 16'b0000001010100000;
            15'd4643: log10_cal = 16'b0000001010100000;
            15'd4644: log10_cal = 16'b0000001010100000;
            15'd4645: log10_cal = 16'b0000001010100000;
            15'd4646: log10_cal = 16'b0000001010100000;
            15'd4647: log10_cal = 16'b0000001010100000;
            15'd4648: log10_cal = 16'b0000001010100000;
            15'd4649: log10_cal = 16'b0000001010100000;
            15'd4650: log10_cal = 16'b0000001010100000;
            15'd4651: log10_cal = 16'b0000001010100001;
            15'd4652: log10_cal = 16'b0000001010100001;
            15'd4653: log10_cal = 16'b0000001010100001;
            15'd4654: log10_cal = 16'b0000001010100001;
            15'd4655: log10_cal = 16'b0000001010100001;
            15'd4656: log10_cal = 16'b0000001010100001;
            15'd4657: log10_cal = 16'b0000001010100001;
            15'd4658: log10_cal = 16'b0000001010100001;
            15'd4659: log10_cal = 16'b0000001010100001;
            15'd4660: log10_cal = 16'b0000001010100001;
            15'd4661: log10_cal = 16'b0000001010100001;
            15'd4662: log10_cal = 16'b0000001010100010;
            15'd4663: log10_cal = 16'b0000001010100010;
            15'd4664: log10_cal = 16'b0000001010100010;
            15'd4665: log10_cal = 16'b0000001010100010;
            15'd4666: log10_cal = 16'b0000001010100010;
            15'd4667: log10_cal = 16'b0000001010100010;
            15'd4668: log10_cal = 16'b0000001010100010;
            15'd4669: log10_cal = 16'b0000001010100010;
            15'd4670: log10_cal = 16'b0000001010100010;
            15'd4671: log10_cal = 16'b0000001010100010;
            15'd4672: log10_cal = 16'b0000001010100011;
            15'd4673: log10_cal = 16'b0000001010100011;
            15'd4674: log10_cal = 16'b0000001010100011;
            15'd4675: log10_cal = 16'b0000001010100011;
            15'd4676: log10_cal = 16'b0000001010100011;
            15'd4677: log10_cal = 16'b0000001010100011;
            15'd4678: log10_cal = 16'b0000001010100011;
            15'd4679: log10_cal = 16'b0000001010100011;
            15'd4680: log10_cal = 16'b0000001010100011;
            15'd4681: log10_cal = 16'b0000001010100011;
            15'd4682: log10_cal = 16'b0000001010100011;
            15'd4683: log10_cal = 16'b0000001010100100;
            15'd4684: log10_cal = 16'b0000001010100100;
            15'd4685: log10_cal = 16'b0000001010100100;
            15'd4686: log10_cal = 16'b0000001010100100;
            15'd4687: log10_cal = 16'b0000001010100100;
            15'd4688: log10_cal = 16'b0000001010100100;
            15'd4689: log10_cal = 16'b0000001010100100;
            15'd4690: log10_cal = 16'b0000001010100100;
            15'd4691: log10_cal = 16'b0000001010100100;
            15'd4692: log10_cal = 16'b0000001010100100;
            15'd4693: log10_cal = 16'b0000001010100101;
            15'd4694: log10_cal = 16'b0000001010100101;
            15'd4695: log10_cal = 16'b0000001010100101;
            15'd4696: log10_cal = 16'b0000001010100101;
            15'd4697: log10_cal = 16'b0000001010100101;
            15'd4698: log10_cal = 16'b0000001010100101;
            15'd4699: log10_cal = 16'b0000001010100101;
            15'd4700: log10_cal = 16'b0000001010100101;
            15'd4701: log10_cal = 16'b0000001010100101;
            15'd4702: log10_cal = 16'b0000001010100101;
            15'd4703: log10_cal = 16'b0000001010100101;
            15'd4704: log10_cal = 16'b0000001010100110;
            15'd4705: log10_cal = 16'b0000001010100110;
            15'd4706: log10_cal = 16'b0000001010100110;
            15'd4707: log10_cal = 16'b0000001010100110;
            15'd4708: log10_cal = 16'b0000001010100110;
            15'd4709: log10_cal = 16'b0000001010100110;
            15'd4710: log10_cal = 16'b0000001010100110;
            15'd4711: log10_cal = 16'b0000001010100110;
            15'd4712: log10_cal = 16'b0000001010100110;
            15'd4713: log10_cal = 16'b0000001010100110;
            15'd4714: log10_cal = 16'b0000001010100111;
            15'd4715: log10_cal = 16'b0000001010100111;
            15'd4716: log10_cal = 16'b0000001010100111;
            15'd4717: log10_cal = 16'b0000001010100111;
            15'd4718: log10_cal = 16'b0000001010100111;
            15'd4719: log10_cal = 16'b0000001010100111;
            15'd4720: log10_cal = 16'b0000001010100111;
            15'd4721: log10_cal = 16'b0000001010100111;
            15'd4722: log10_cal = 16'b0000001010100111;
            15'd4723: log10_cal = 16'b0000001010100111;
            15'd4724: log10_cal = 16'b0000001010100111;
            15'd4725: log10_cal = 16'b0000001010101000;
            15'd4726: log10_cal = 16'b0000001010101000;
            15'd4727: log10_cal = 16'b0000001010101000;
            15'd4728: log10_cal = 16'b0000001010101000;
            15'd4729: log10_cal = 16'b0000001010101000;
            15'd4730: log10_cal = 16'b0000001010101000;
            15'd4731: log10_cal = 16'b0000001010101000;
            15'd4732: log10_cal = 16'b0000001010101000;
            15'd4733: log10_cal = 16'b0000001010101000;
            15'd4734: log10_cal = 16'b0000001010101000;
            15'd4735: log10_cal = 16'b0000001010101000;
            15'd4736: log10_cal = 16'b0000001010101001;
            15'd4737: log10_cal = 16'b0000001010101001;
            15'd4738: log10_cal = 16'b0000001010101001;
            15'd4739: log10_cal = 16'b0000001010101001;
            15'd4740: log10_cal = 16'b0000001010101001;
            15'd4741: log10_cal = 16'b0000001010101001;
            15'd4742: log10_cal = 16'b0000001010101001;
            15'd4743: log10_cal = 16'b0000001010101001;
            15'd4744: log10_cal = 16'b0000001010101001;
            15'd4745: log10_cal = 16'b0000001010101001;
            15'd4746: log10_cal = 16'b0000001010101010;
            15'd4747: log10_cal = 16'b0000001010101010;
            15'd4748: log10_cal = 16'b0000001010101010;
            15'd4749: log10_cal = 16'b0000001010101010;
            15'd4750: log10_cal = 16'b0000001010101010;
            15'd4751: log10_cal = 16'b0000001010101010;
            15'd4752: log10_cal = 16'b0000001010101010;
            15'd4753: log10_cal = 16'b0000001010101010;
            15'd4754: log10_cal = 16'b0000001010101010;
            15'd4755: log10_cal = 16'b0000001010101010;
            15'd4756: log10_cal = 16'b0000001010101010;
            15'd4757: log10_cal = 16'b0000001010101011;
            15'd4758: log10_cal = 16'b0000001010101011;
            15'd4759: log10_cal = 16'b0000001010101011;
            15'd4760: log10_cal = 16'b0000001010101011;
            15'd4761: log10_cal = 16'b0000001010101011;
            15'd4762: log10_cal = 16'b0000001010101011;
            15'd4763: log10_cal = 16'b0000001010101011;
            15'd4764: log10_cal = 16'b0000001010101011;
            15'd4765: log10_cal = 16'b0000001010101011;
            15'd4766: log10_cal = 16'b0000001010101011;
            15'd4767: log10_cal = 16'b0000001010101011;
            15'd4768: log10_cal = 16'b0000001010101100;
            15'd4769: log10_cal = 16'b0000001010101100;
            15'd4770: log10_cal = 16'b0000001010101100;
            15'd4771: log10_cal = 16'b0000001010101100;
            15'd4772: log10_cal = 16'b0000001010101100;
            15'd4773: log10_cal = 16'b0000001010101100;
            15'd4774: log10_cal = 16'b0000001010101100;
            15'd4775: log10_cal = 16'b0000001010101100;
            15'd4776: log10_cal = 16'b0000001010101100;
            15'd4777: log10_cal = 16'b0000001010101100;
            15'd4778: log10_cal = 16'b0000001010101101;
            15'd4779: log10_cal = 16'b0000001010101101;
            15'd4780: log10_cal = 16'b0000001010101101;
            15'd4781: log10_cal = 16'b0000001010101101;
            15'd4782: log10_cal = 16'b0000001010101101;
            15'd4783: log10_cal = 16'b0000001010101101;
            15'd4784: log10_cal = 16'b0000001010101101;
            15'd4785: log10_cal = 16'b0000001010101101;
            15'd4786: log10_cal = 16'b0000001010101101;
            15'd4787: log10_cal = 16'b0000001010101101;
            15'd4788: log10_cal = 16'b0000001010101101;
            15'd4789: log10_cal = 16'b0000001010101110;
            15'd4790: log10_cal = 16'b0000001010101110;
            15'd4791: log10_cal = 16'b0000001010101110;
            15'd4792: log10_cal = 16'b0000001010101110;
            15'd4793: log10_cal = 16'b0000001010101110;
            15'd4794: log10_cal = 16'b0000001010101110;
            15'd4795: log10_cal = 16'b0000001010101110;
            15'd4796: log10_cal = 16'b0000001010101110;
            15'd4797: log10_cal = 16'b0000001010101110;
            15'd4798: log10_cal = 16'b0000001010101110;
            15'd4799: log10_cal = 16'b0000001010101110;
            15'd4800: log10_cal = 16'b0000001010101111;
            15'd4801: log10_cal = 16'b0000001010101111;
            15'd4802: log10_cal = 16'b0000001010101111;
            15'd4803: log10_cal = 16'b0000001010101111;
            15'd4804: log10_cal = 16'b0000001010101111;
            15'd4805: log10_cal = 16'b0000001010101111;
            15'd4806: log10_cal = 16'b0000001010101111;
            15'd4807: log10_cal = 16'b0000001010101111;
            15'd4808: log10_cal = 16'b0000001010101111;
            15'd4809: log10_cal = 16'b0000001010101111;
            15'd4810: log10_cal = 16'b0000001010101111;
            15'd4811: log10_cal = 16'b0000001010110000;
            15'd4812: log10_cal = 16'b0000001010110000;
            15'd4813: log10_cal = 16'b0000001010110000;
            15'd4814: log10_cal = 16'b0000001010110000;
            15'd4815: log10_cal = 16'b0000001010110000;
            15'd4816: log10_cal = 16'b0000001010110000;
            15'd4817: log10_cal = 16'b0000001010110000;
            15'd4818: log10_cal = 16'b0000001010110000;
            15'd4819: log10_cal = 16'b0000001010110000;
            15'd4820: log10_cal = 16'b0000001010110000;
            15'd4821: log10_cal = 16'b0000001010110000;
            15'd4822: log10_cal = 16'b0000001010110001;
            15'd4823: log10_cal = 16'b0000001010110001;
            15'd4824: log10_cal = 16'b0000001010110001;
            15'd4825: log10_cal = 16'b0000001010110001;
            15'd4826: log10_cal = 16'b0000001010110001;
            15'd4827: log10_cal = 16'b0000001010110001;
            15'd4828: log10_cal = 16'b0000001010110001;
            15'd4829: log10_cal = 16'b0000001010110001;
            15'd4830: log10_cal = 16'b0000001010110001;
            15'd4831: log10_cal = 16'b0000001010110001;
            15'd4832: log10_cal = 16'b0000001010110001;
            15'd4833: log10_cal = 16'b0000001010110010;
            15'd4834: log10_cal = 16'b0000001010110010;
            15'd4835: log10_cal = 16'b0000001010110010;
            15'd4836: log10_cal = 16'b0000001010110010;
            15'd4837: log10_cal = 16'b0000001010110010;
            15'd4838: log10_cal = 16'b0000001010110010;
            15'd4839: log10_cal = 16'b0000001010110010;
            15'd4840: log10_cal = 16'b0000001010110010;
            15'd4841: log10_cal = 16'b0000001010110010;
            15'd4842: log10_cal = 16'b0000001010110010;
            15'd4843: log10_cal = 16'b0000001010110011;
            15'd4844: log10_cal = 16'b0000001010110011;
            15'd4845: log10_cal = 16'b0000001010110011;
            15'd4846: log10_cal = 16'b0000001010110011;
            15'd4847: log10_cal = 16'b0000001010110011;
            15'd4848: log10_cal = 16'b0000001010110011;
            15'd4849: log10_cal = 16'b0000001010110011;
            15'd4850: log10_cal = 16'b0000001010110011;
            15'd4851: log10_cal = 16'b0000001010110011;
            15'd4852: log10_cal = 16'b0000001010110011;
            15'd4853: log10_cal = 16'b0000001010110011;
            15'd4854: log10_cal = 16'b0000001010110100;
            15'd4855: log10_cal = 16'b0000001010110100;
            15'd4856: log10_cal = 16'b0000001010110100;
            15'd4857: log10_cal = 16'b0000001010110100;
            15'd4858: log10_cal = 16'b0000001010110100;
            15'd4859: log10_cal = 16'b0000001010110100;
            15'd4860: log10_cal = 16'b0000001010110100;
            15'd4861: log10_cal = 16'b0000001010110100;
            15'd4862: log10_cal = 16'b0000001010110100;
            15'd4863: log10_cal = 16'b0000001010110100;
            15'd4864: log10_cal = 16'b0000001010110100;
            15'd4865: log10_cal = 16'b0000001010110101;
            15'd4866: log10_cal = 16'b0000001010110101;
            15'd4867: log10_cal = 16'b0000001010110101;
            15'd4868: log10_cal = 16'b0000001010110101;
            15'd4869: log10_cal = 16'b0000001010110101;
            15'd4870: log10_cal = 16'b0000001010110101;
            15'd4871: log10_cal = 16'b0000001010110101;
            15'd4872: log10_cal = 16'b0000001010110101;
            15'd4873: log10_cal = 16'b0000001010110101;
            15'd4874: log10_cal = 16'b0000001010110101;
            15'd4875: log10_cal = 16'b0000001010110101;
            15'd4876: log10_cal = 16'b0000001010110110;
            15'd4877: log10_cal = 16'b0000001010110110;
            15'd4878: log10_cal = 16'b0000001010110110;
            15'd4879: log10_cal = 16'b0000001010110110;
            15'd4880: log10_cal = 16'b0000001010110110;
            15'd4881: log10_cal = 16'b0000001010110110;
            15'd4882: log10_cal = 16'b0000001010110110;
            15'd4883: log10_cal = 16'b0000001010110110;
            15'd4884: log10_cal = 16'b0000001010110110;
            15'd4885: log10_cal = 16'b0000001010110110;
            15'd4886: log10_cal = 16'b0000001010110110;
            15'd4887: log10_cal = 16'b0000001010110111;
            15'd4888: log10_cal = 16'b0000001010110111;
            15'd4889: log10_cal = 16'b0000001010110111;
            15'd4890: log10_cal = 16'b0000001010110111;
            15'd4891: log10_cal = 16'b0000001010110111;
            15'd4892: log10_cal = 16'b0000001010110111;
            15'd4893: log10_cal = 16'b0000001010110111;
            15'd4894: log10_cal = 16'b0000001010110111;
            15'd4895: log10_cal = 16'b0000001010110111;
            15'd4896: log10_cal = 16'b0000001010110111;
            15'd4897: log10_cal = 16'b0000001010110111;
            15'd4898: log10_cal = 16'b0000001010111000;
            15'd4899: log10_cal = 16'b0000001010111000;
            15'd4900: log10_cal = 16'b0000001010111000;
            15'd4901: log10_cal = 16'b0000001010111000;
            15'd4902: log10_cal = 16'b0000001010111000;
            15'd4903: log10_cal = 16'b0000001010111000;
            15'd4904: log10_cal = 16'b0000001010111000;
            15'd4905: log10_cal = 16'b0000001010111000;
            15'd4906: log10_cal = 16'b0000001010111000;
            15'd4907: log10_cal = 16'b0000001010111000;
            15'd4908: log10_cal = 16'b0000001010111000;
            15'd4909: log10_cal = 16'b0000001010111001;
            15'd4910: log10_cal = 16'b0000001010111001;
            15'd4911: log10_cal = 16'b0000001010111001;
            15'd4912: log10_cal = 16'b0000001010111001;
            15'd4913: log10_cal = 16'b0000001010111001;
            15'd4914: log10_cal = 16'b0000001010111001;
            15'd4915: log10_cal = 16'b0000001010111001;
            15'd4916: log10_cal = 16'b0000001010111001;
            15'd4917: log10_cal = 16'b0000001010111001;
            15'd4918: log10_cal = 16'b0000001010111001;
            15'd4919: log10_cal = 16'b0000001010111001;
            15'd4920: log10_cal = 16'b0000001010111010;
            15'd4921: log10_cal = 16'b0000001010111010;
            15'd4922: log10_cal = 16'b0000001010111010;
            15'd4923: log10_cal = 16'b0000001010111010;
            15'd4924: log10_cal = 16'b0000001010111010;
            15'd4925: log10_cal = 16'b0000001010111010;
            15'd4926: log10_cal = 16'b0000001010111010;
            15'd4927: log10_cal = 16'b0000001010111010;
            15'd4928: log10_cal = 16'b0000001010111010;
            15'd4929: log10_cal = 16'b0000001010111010;
            15'd4930: log10_cal = 16'b0000001010111010;
            15'd4931: log10_cal = 16'b0000001010111011;
            15'd4932: log10_cal = 16'b0000001010111011;
            15'd4933: log10_cal = 16'b0000001010111011;
            15'd4934: log10_cal = 16'b0000001010111011;
            15'd4935: log10_cal = 16'b0000001010111011;
            15'd4936: log10_cal = 16'b0000001010111011;
            15'd4937: log10_cal = 16'b0000001010111011;
            15'd4938: log10_cal = 16'b0000001010111011;
            15'd4939: log10_cal = 16'b0000001010111011;
            15'd4940: log10_cal = 16'b0000001010111011;
            15'd4941: log10_cal = 16'b0000001010111011;
            15'd4942: log10_cal = 16'b0000001010111100;
            15'd4943: log10_cal = 16'b0000001010111100;
            15'd4944: log10_cal = 16'b0000001010111100;
            15'd4945: log10_cal = 16'b0000001010111100;
            15'd4946: log10_cal = 16'b0000001010111100;
            15'd4947: log10_cal = 16'b0000001010111100;
            15'd4948: log10_cal = 16'b0000001010111100;
            15'd4949: log10_cal = 16'b0000001010111100;
            15'd4950: log10_cal = 16'b0000001010111100;
            15'd4951: log10_cal = 16'b0000001010111100;
            15'd4952: log10_cal = 16'b0000001010111100;
            15'd4953: log10_cal = 16'b0000001010111100;
            15'd4954: log10_cal = 16'b0000001010111101;
            15'd4955: log10_cal = 16'b0000001010111101;
            15'd4956: log10_cal = 16'b0000001010111101;
            15'd4957: log10_cal = 16'b0000001010111101;
            15'd4958: log10_cal = 16'b0000001010111101;
            15'd4959: log10_cal = 16'b0000001010111101;
            15'd4960: log10_cal = 16'b0000001010111101;
            15'd4961: log10_cal = 16'b0000001010111101;
            15'd4962: log10_cal = 16'b0000001010111101;
            15'd4963: log10_cal = 16'b0000001010111101;
            15'd4964: log10_cal = 16'b0000001010111101;
            15'd4965: log10_cal = 16'b0000001010111110;
            15'd4966: log10_cal = 16'b0000001010111110;
            15'd4967: log10_cal = 16'b0000001010111110;
            15'd4968: log10_cal = 16'b0000001010111110;
            15'd4969: log10_cal = 16'b0000001010111110;
            15'd4970: log10_cal = 16'b0000001010111110;
            15'd4971: log10_cal = 16'b0000001010111110;
            15'd4972: log10_cal = 16'b0000001010111110;
            15'd4973: log10_cal = 16'b0000001010111110;
            15'd4974: log10_cal = 16'b0000001010111110;
            15'd4975: log10_cal = 16'b0000001010111110;
            15'd4976: log10_cal = 16'b0000001010111111;
            15'd4977: log10_cal = 16'b0000001010111111;
            15'd4978: log10_cal = 16'b0000001010111111;
            15'd4979: log10_cal = 16'b0000001010111111;
            15'd4980: log10_cal = 16'b0000001010111111;
            15'd4981: log10_cal = 16'b0000001010111111;
            15'd4982: log10_cal = 16'b0000001010111111;
            15'd4983: log10_cal = 16'b0000001010111111;
            15'd4984: log10_cal = 16'b0000001010111111;
            15'd4985: log10_cal = 16'b0000001010111111;
            15'd4986: log10_cal = 16'b0000001010111111;
            15'd4987: log10_cal = 16'b0000001011000000;
            15'd4988: log10_cal = 16'b0000001011000000;
            15'd4989: log10_cal = 16'b0000001011000000;
            15'd4990: log10_cal = 16'b0000001011000000;
            15'd4991: log10_cal = 16'b0000001011000000;
            15'd4992: log10_cal = 16'b0000001011000000;
            15'd4993: log10_cal = 16'b0000001011000000;
            15'd4994: log10_cal = 16'b0000001011000000;
            15'd4995: log10_cal = 16'b0000001011000000;
            15'd4996: log10_cal = 16'b0000001011000000;
            15'd4997: log10_cal = 16'b0000001011000000;
            15'd4998: log10_cal = 16'b0000001011000001;
            15'd4999: log10_cal = 16'b0000001011000001;
            15'd5000: log10_cal = 16'b0000001011000001;
            15'd5001: log10_cal = 16'b0000001011000001;
            15'd5002: log10_cal = 16'b0000001011000001;
            15'd5003: log10_cal = 16'b0000001011000001;
            15'd5004: log10_cal = 16'b0000001011000001;
            15'd5005: log10_cal = 16'b0000001011000001;
            15'd5006: log10_cal = 16'b0000001011000001;
            15'd5007: log10_cal = 16'b0000001011000001;
            15'd5008: log10_cal = 16'b0000001011000001;
            15'd5009: log10_cal = 16'b0000001011000001;
            15'd5010: log10_cal = 16'b0000001011000010;
            15'd5011: log10_cal = 16'b0000001011000010;
            15'd5012: log10_cal = 16'b0000001011000010;
            15'd5013: log10_cal = 16'b0000001011000010;
            15'd5014: log10_cal = 16'b0000001011000010;
            15'd5015: log10_cal = 16'b0000001011000010;
            15'd5016: log10_cal = 16'b0000001011000010;
            15'd5017: log10_cal = 16'b0000001011000010;
            15'd5018: log10_cal = 16'b0000001011000010;
            15'd5019: log10_cal = 16'b0000001011000010;
            15'd5020: log10_cal = 16'b0000001011000010;
            15'd5021: log10_cal = 16'b0000001011000011;
            15'd5022: log10_cal = 16'b0000001011000011;
            15'd5023: log10_cal = 16'b0000001011000011;
            15'd5024: log10_cal = 16'b0000001011000011;
            15'd5025: log10_cal = 16'b0000001011000011;
            15'd5026: log10_cal = 16'b0000001011000011;
            15'd5027: log10_cal = 16'b0000001011000011;
            15'd5028: log10_cal = 16'b0000001011000011;
            15'd5029: log10_cal = 16'b0000001011000011;
            15'd5030: log10_cal = 16'b0000001011000011;
            15'd5031: log10_cal = 16'b0000001011000011;
            15'd5032: log10_cal = 16'b0000001011000100;
            15'd5033: log10_cal = 16'b0000001011000100;
            15'd5034: log10_cal = 16'b0000001011000100;
            15'd5035: log10_cal = 16'b0000001011000100;
            15'd5036: log10_cal = 16'b0000001011000100;
            15'd5037: log10_cal = 16'b0000001011000100;
            15'd5038: log10_cal = 16'b0000001011000100;
            15'd5039: log10_cal = 16'b0000001011000100;
            15'd5040: log10_cal = 16'b0000001011000100;
            15'd5041: log10_cal = 16'b0000001011000100;
            15'd5042: log10_cal = 16'b0000001011000100;
            15'd5043: log10_cal = 16'b0000001011000101;
            15'd5044: log10_cal = 16'b0000001011000101;
            15'd5045: log10_cal = 16'b0000001011000101;
            15'd5046: log10_cal = 16'b0000001011000101;
            15'd5047: log10_cal = 16'b0000001011000101;
            15'd5048: log10_cal = 16'b0000001011000101;
            15'd5049: log10_cal = 16'b0000001011000101;
            15'd5050: log10_cal = 16'b0000001011000101;
            15'd5051: log10_cal = 16'b0000001011000101;
            15'd5052: log10_cal = 16'b0000001011000101;
            15'd5053: log10_cal = 16'b0000001011000101;
            15'd5054: log10_cal = 16'b0000001011000101;
            15'd5055: log10_cal = 16'b0000001011000110;
            15'd5056: log10_cal = 16'b0000001011000110;
            15'd5057: log10_cal = 16'b0000001011000110;
            15'd5058: log10_cal = 16'b0000001011000110;
            15'd5059: log10_cal = 16'b0000001011000110;
            15'd5060: log10_cal = 16'b0000001011000110;
            15'd5061: log10_cal = 16'b0000001011000110;
            15'd5062: log10_cal = 16'b0000001011000110;
            15'd5063: log10_cal = 16'b0000001011000110;
            15'd5064: log10_cal = 16'b0000001011000110;
            15'd5065: log10_cal = 16'b0000001011000110;
            15'd5066: log10_cal = 16'b0000001011000111;
            15'd5067: log10_cal = 16'b0000001011000111;
            15'd5068: log10_cal = 16'b0000001011000111;
            15'd5069: log10_cal = 16'b0000001011000111;
            15'd5070: log10_cal = 16'b0000001011000111;
            15'd5071: log10_cal = 16'b0000001011000111;
            15'd5072: log10_cal = 16'b0000001011000111;
            15'd5073: log10_cal = 16'b0000001011000111;
            15'd5074: log10_cal = 16'b0000001011000111;
            15'd5075: log10_cal = 16'b0000001011000111;
            15'd5076: log10_cal = 16'b0000001011000111;
            15'd5077: log10_cal = 16'b0000001011000111;
            15'd5078: log10_cal = 16'b0000001011001000;
            15'd5079: log10_cal = 16'b0000001011001000;
            15'd5080: log10_cal = 16'b0000001011001000;
            15'd5081: log10_cal = 16'b0000001011001000;
            15'd5082: log10_cal = 16'b0000001011001000;
            15'd5083: log10_cal = 16'b0000001011001000;
            15'd5084: log10_cal = 16'b0000001011001000;
            15'd5085: log10_cal = 16'b0000001011001000;
            15'd5086: log10_cal = 16'b0000001011001000;
            15'd5087: log10_cal = 16'b0000001011001000;
            15'd5088: log10_cal = 16'b0000001011001000;
            15'd5089: log10_cal = 16'b0000001011001001;
            15'd5090: log10_cal = 16'b0000001011001001;
            15'd5091: log10_cal = 16'b0000001011001001;
            15'd5092: log10_cal = 16'b0000001011001001;
            15'd5093: log10_cal = 16'b0000001011001001;
            15'd5094: log10_cal = 16'b0000001011001001;
            15'd5095: log10_cal = 16'b0000001011001001;
            15'd5096: log10_cal = 16'b0000001011001001;
            15'd5097: log10_cal = 16'b0000001011001001;
            15'd5098: log10_cal = 16'b0000001011001001;
            15'd5099: log10_cal = 16'b0000001011001001;
            15'd5100: log10_cal = 16'b0000001011001010;
            15'd5101: log10_cal = 16'b0000001011001010;
            15'd5102: log10_cal = 16'b0000001011001010;
            15'd5103: log10_cal = 16'b0000001011001010;
            15'd5104: log10_cal = 16'b0000001011001010;
            15'd5105: log10_cal = 16'b0000001011001010;
            15'd5106: log10_cal = 16'b0000001011001010;
            15'd5107: log10_cal = 16'b0000001011001010;
            15'd5108: log10_cal = 16'b0000001011001010;
            15'd5109: log10_cal = 16'b0000001011001010;
            15'd5110: log10_cal = 16'b0000001011001010;
            15'd5111: log10_cal = 16'b0000001011001010;
            15'd5112: log10_cal = 16'b0000001011001011;
            15'd5113: log10_cal = 16'b0000001011001011;
            15'd5114: log10_cal = 16'b0000001011001011;
            15'd5115: log10_cal = 16'b0000001011001011;
            15'd5116: log10_cal = 16'b0000001011001011;
            15'd5117: log10_cal = 16'b0000001011001011;
            15'd5118: log10_cal = 16'b0000001011001011;
            15'd5119: log10_cal = 16'b0000001011001011;
            15'd5120: log10_cal = 16'b0000001011001011;
            15'd5121: log10_cal = 16'b0000001011001011;
            15'd5122: log10_cal = 16'b0000001011001011;
            15'd5123: log10_cal = 16'b0000001011001100;
            15'd5124: log10_cal = 16'b0000001011001100;
            15'd5125: log10_cal = 16'b0000001011001100;
            15'd5126: log10_cal = 16'b0000001011001100;
            15'd5127: log10_cal = 16'b0000001011001100;
            15'd5128: log10_cal = 16'b0000001011001100;
            15'd5129: log10_cal = 16'b0000001011001100;
            15'd5130: log10_cal = 16'b0000001011001100;
            15'd5131: log10_cal = 16'b0000001011001100;
            15'd5132: log10_cal = 16'b0000001011001100;
            15'd5133: log10_cal = 16'b0000001011001100;
            15'd5134: log10_cal = 16'b0000001011001100;
            15'd5135: log10_cal = 16'b0000001011001101;
            15'd5136: log10_cal = 16'b0000001011001101;
            15'd5137: log10_cal = 16'b0000001011001101;
            15'd5138: log10_cal = 16'b0000001011001101;
            15'd5139: log10_cal = 16'b0000001011001101;
            15'd5140: log10_cal = 16'b0000001011001101;
            15'd5141: log10_cal = 16'b0000001011001101;
            15'd5142: log10_cal = 16'b0000001011001101;
            15'd5143: log10_cal = 16'b0000001011001101;
            15'd5144: log10_cal = 16'b0000001011001101;
            15'd5145: log10_cal = 16'b0000001011001101;
            15'd5146: log10_cal = 16'b0000001011001101;
            15'd5147: log10_cal = 16'b0000001011001110;
            15'd5148: log10_cal = 16'b0000001011001110;
            15'd5149: log10_cal = 16'b0000001011001110;
            15'd5150: log10_cal = 16'b0000001011001110;
            15'd5151: log10_cal = 16'b0000001011001110;
            15'd5152: log10_cal = 16'b0000001011001110;
            15'd5153: log10_cal = 16'b0000001011001110;
            15'd5154: log10_cal = 16'b0000001011001110;
            15'd5155: log10_cal = 16'b0000001011001110;
            15'd5156: log10_cal = 16'b0000001011001110;
            15'd5157: log10_cal = 16'b0000001011001110;
            15'd5158: log10_cal = 16'b0000001011001111;
            15'd5159: log10_cal = 16'b0000001011001111;
            15'd5160: log10_cal = 16'b0000001011001111;
            15'd5161: log10_cal = 16'b0000001011001111;
            15'd5162: log10_cal = 16'b0000001011001111;
            15'd5163: log10_cal = 16'b0000001011001111;
            15'd5164: log10_cal = 16'b0000001011001111;
            15'd5165: log10_cal = 16'b0000001011001111;
            15'd5166: log10_cal = 16'b0000001011001111;
            15'd5167: log10_cal = 16'b0000001011001111;
            15'd5168: log10_cal = 16'b0000001011001111;
            15'd5169: log10_cal = 16'b0000001011001111;
            15'd5170: log10_cal = 16'b0000001011010000;
            15'd5171: log10_cal = 16'b0000001011010000;
            15'd5172: log10_cal = 16'b0000001011010000;
            15'd5173: log10_cal = 16'b0000001011010000;
            15'd5174: log10_cal = 16'b0000001011010000;
            15'd5175: log10_cal = 16'b0000001011010000;
            15'd5176: log10_cal = 16'b0000001011010000;
            15'd5177: log10_cal = 16'b0000001011010000;
            15'd5178: log10_cal = 16'b0000001011010000;
            15'd5179: log10_cal = 16'b0000001011010000;
            15'd5180: log10_cal = 16'b0000001011010000;
            15'd5181: log10_cal = 16'b0000001011010001;
            15'd5182: log10_cal = 16'b0000001011010001;
            15'd5183: log10_cal = 16'b0000001011010001;
            15'd5184: log10_cal = 16'b0000001011010001;
            15'd5185: log10_cal = 16'b0000001011010001;
            15'd5186: log10_cal = 16'b0000001011010001;
            15'd5187: log10_cal = 16'b0000001011010001;
            15'd5188: log10_cal = 16'b0000001011010001;
            15'd5189: log10_cal = 16'b0000001011010001;
            15'd5190: log10_cal = 16'b0000001011010001;
            15'd5191: log10_cal = 16'b0000001011010001;
            15'd5192: log10_cal = 16'b0000001011010001;
            15'd5193: log10_cal = 16'b0000001011010010;
            15'd5194: log10_cal = 16'b0000001011010010;
            15'd5195: log10_cal = 16'b0000001011010010;
            15'd5196: log10_cal = 16'b0000001011010010;
            15'd5197: log10_cal = 16'b0000001011010010;
            15'd5198: log10_cal = 16'b0000001011010010;
            15'd5199: log10_cal = 16'b0000001011010010;
            15'd5200: log10_cal = 16'b0000001011010010;
            15'd5201: log10_cal = 16'b0000001011010010;
            15'd5202: log10_cal = 16'b0000001011010010;
            15'd5203: log10_cal = 16'b0000001011010010;
            15'd5204: log10_cal = 16'b0000001011010010;
            15'd5205: log10_cal = 16'b0000001011010011;
            15'd5206: log10_cal = 16'b0000001011010011;
            15'd5207: log10_cal = 16'b0000001011010011;
            15'd5208: log10_cal = 16'b0000001011010011;
            15'd5209: log10_cal = 16'b0000001011010011;
            15'd5210: log10_cal = 16'b0000001011010011;
            15'd5211: log10_cal = 16'b0000001011010011;
            15'd5212: log10_cal = 16'b0000001011010011;
            15'd5213: log10_cal = 16'b0000001011010011;
            15'd5214: log10_cal = 16'b0000001011010011;
            15'd5215: log10_cal = 16'b0000001011010011;
            15'd5216: log10_cal = 16'b0000001011010100;
            15'd5217: log10_cal = 16'b0000001011010100;
            15'd5218: log10_cal = 16'b0000001011010100;
            15'd5219: log10_cal = 16'b0000001011010100;
            15'd5220: log10_cal = 16'b0000001011010100;
            15'd5221: log10_cal = 16'b0000001011010100;
            15'd5222: log10_cal = 16'b0000001011010100;
            15'd5223: log10_cal = 16'b0000001011010100;
            15'd5224: log10_cal = 16'b0000001011010100;
            15'd5225: log10_cal = 16'b0000001011010100;
            15'd5226: log10_cal = 16'b0000001011010100;
            15'd5227: log10_cal = 16'b0000001011010100;
            15'd5228: log10_cal = 16'b0000001011010101;
            15'd5229: log10_cal = 16'b0000001011010101;
            15'd5230: log10_cal = 16'b0000001011010101;
            15'd5231: log10_cal = 16'b0000001011010101;
            15'd5232: log10_cal = 16'b0000001011010101;
            15'd5233: log10_cal = 16'b0000001011010101;
            15'd5234: log10_cal = 16'b0000001011010101;
            15'd5235: log10_cal = 16'b0000001011010101;
            15'd5236: log10_cal = 16'b0000001011010101;
            15'd5237: log10_cal = 16'b0000001011010101;
            15'd5238: log10_cal = 16'b0000001011010101;
            15'd5239: log10_cal = 16'b0000001011010101;
            15'd5240: log10_cal = 16'b0000001011010110;
            15'd5241: log10_cal = 16'b0000001011010110;
            15'd5242: log10_cal = 16'b0000001011010110;
            15'd5243: log10_cal = 16'b0000001011010110;
            15'd5244: log10_cal = 16'b0000001011010110;
            15'd5245: log10_cal = 16'b0000001011010110;
            15'd5246: log10_cal = 16'b0000001011010110;
            15'd5247: log10_cal = 16'b0000001011010110;
            15'd5248: log10_cal = 16'b0000001011010110;
            15'd5249: log10_cal = 16'b0000001011010110;
            15'd5250: log10_cal = 16'b0000001011010110;
            15'd5251: log10_cal = 16'b0000001011010110;
            15'd5252: log10_cal = 16'b0000001011010111;
            15'd5253: log10_cal = 16'b0000001011010111;
            15'd5254: log10_cal = 16'b0000001011010111;
            15'd5255: log10_cal = 16'b0000001011010111;
            15'd5256: log10_cal = 16'b0000001011010111;
            15'd5257: log10_cal = 16'b0000001011010111;
            15'd5258: log10_cal = 16'b0000001011010111;
            15'd5259: log10_cal = 16'b0000001011010111;
            15'd5260: log10_cal = 16'b0000001011010111;
            15'd5261: log10_cal = 16'b0000001011010111;
            15'd5262: log10_cal = 16'b0000001011010111;
            15'd5263: log10_cal = 16'b0000001011010111;
            15'd5264: log10_cal = 16'b0000001011011000;
            15'd5265: log10_cal = 16'b0000001011011000;
            15'd5266: log10_cal = 16'b0000001011011000;
            15'd5267: log10_cal = 16'b0000001011011000;
            15'd5268: log10_cal = 16'b0000001011011000;
            15'd5269: log10_cal = 16'b0000001011011000;
            15'd5270: log10_cal = 16'b0000001011011000;
            15'd5271: log10_cal = 16'b0000001011011000;
            15'd5272: log10_cal = 16'b0000001011011000;
            15'd5273: log10_cal = 16'b0000001011011000;
            15'd5274: log10_cal = 16'b0000001011011000;
            15'd5275: log10_cal = 16'b0000001011011001;
            15'd5276: log10_cal = 16'b0000001011011001;
            15'd5277: log10_cal = 16'b0000001011011001;
            15'd5278: log10_cal = 16'b0000001011011001;
            15'd5279: log10_cal = 16'b0000001011011001;
            15'd5280: log10_cal = 16'b0000001011011001;
            15'd5281: log10_cal = 16'b0000001011011001;
            15'd5282: log10_cal = 16'b0000001011011001;
            15'd5283: log10_cal = 16'b0000001011011001;
            15'd5284: log10_cal = 16'b0000001011011001;
            15'd5285: log10_cal = 16'b0000001011011001;
            15'd5286: log10_cal = 16'b0000001011011001;
            15'd5287: log10_cal = 16'b0000001011011010;
            15'd5288: log10_cal = 16'b0000001011011010;
            15'd5289: log10_cal = 16'b0000001011011010;
            15'd5290: log10_cal = 16'b0000001011011010;
            15'd5291: log10_cal = 16'b0000001011011010;
            15'd5292: log10_cal = 16'b0000001011011010;
            15'd5293: log10_cal = 16'b0000001011011010;
            15'd5294: log10_cal = 16'b0000001011011010;
            15'd5295: log10_cal = 16'b0000001011011010;
            15'd5296: log10_cal = 16'b0000001011011010;
            15'd5297: log10_cal = 16'b0000001011011010;
            15'd5298: log10_cal = 16'b0000001011011010;
            15'd5299: log10_cal = 16'b0000001011011011;
            15'd5300: log10_cal = 16'b0000001011011011;
            15'd5301: log10_cal = 16'b0000001011011011;
            15'd5302: log10_cal = 16'b0000001011011011;
            15'd5303: log10_cal = 16'b0000001011011011;
            15'd5304: log10_cal = 16'b0000001011011011;
            15'd5305: log10_cal = 16'b0000001011011011;
            15'd5306: log10_cal = 16'b0000001011011011;
            15'd5307: log10_cal = 16'b0000001011011011;
            15'd5308: log10_cal = 16'b0000001011011011;
            15'd5309: log10_cal = 16'b0000001011011011;
            15'd5310: log10_cal = 16'b0000001011011011;
            15'd5311: log10_cal = 16'b0000001011011100;
            15'd5312: log10_cal = 16'b0000001011011100;
            15'd5313: log10_cal = 16'b0000001011011100;
            15'd5314: log10_cal = 16'b0000001011011100;
            15'd5315: log10_cal = 16'b0000001011011100;
            15'd5316: log10_cal = 16'b0000001011011100;
            15'd5317: log10_cal = 16'b0000001011011100;
            15'd5318: log10_cal = 16'b0000001011011100;
            15'd5319: log10_cal = 16'b0000001011011100;
            15'd5320: log10_cal = 16'b0000001011011100;
            15'd5321: log10_cal = 16'b0000001011011100;
            15'd5322: log10_cal = 16'b0000001011011100;
            15'd5323: log10_cal = 16'b0000001011011101;
            15'd5324: log10_cal = 16'b0000001011011101;
            15'd5325: log10_cal = 16'b0000001011011101;
            15'd5326: log10_cal = 16'b0000001011011101;
            15'd5327: log10_cal = 16'b0000001011011101;
            15'd5328: log10_cal = 16'b0000001011011101;
            15'd5329: log10_cal = 16'b0000001011011101;
            15'd5330: log10_cal = 16'b0000001011011101;
            15'd5331: log10_cal = 16'b0000001011011101;
            15'd5332: log10_cal = 16'b0000001011011101;
            15'd5333: log10_cal = 16'b0000001011011101;
            15'd5334: log10_cal = 16'b0000001011011101;
            15'd5335: log10_cal = 16'b0000001011011110;
            15'd5336: log10_cal = 16'b0000001011011110;
            15'd5337: log10_cal = 16'b0000001011011110;
            15'd5338: log10_cal = 16'b0000001011011110;
            15'd5339: log10_cal = 16'b0000001011011110;
            15'd5340: log10_cal = 16'b0000001011011110;
            15'd5341: log10_cal = 16'b0000001011011110;
            15'd5342: log10_cal = 16'b0000001011011110;
            15'd5343: log10_cal = 16'b0000001011011110;
            15'd5344: log10_cal = 16'b0000001011011110;
            15'd5345: log10_cal = 16'b0000001011011110;
            15'd5346: log10_cal = 16'b0000001011011110;
            15'd5347: log10_cal = 16'b0000001011011111;
            15'd5348: log10_cal = 16'b0000001011011111;
            15'd5349: log10_cal = 16'b0000001011011111;
            15'd5350: log10_cal = 16'b0000001011011111;
            15'd5351: log10_cal = 16'b0000001011011111;
            15'd5352: log10_cal = 16'b0000001011011111;
            15'd5353: log10_cal = 16'b0000001011011111;
            15'd5354: log10_cal = 16'b0000001011011111;
            15'd5355: log10_cal = 16'b0000001011011111;
            15'd5356: log10_cal = 16'b0000001011011111;
            15'd5357: log10_cal = 16'b0000001011011111;
            15'd5358: log10_cal = 16'b0000001011011111;
            15'd5359: log10_cal = 16'b0000001011100000;
            15'd5360: log10_cal = 16'b0000001011100000;
            15'd5361: log10_cal = 16'b0000001011100000;
            15'd5362: log10_cal = 16'b0000001011100000;
            15'd5363: log10_cal = 16'b0000001011100000;
            15'd5364: log10_cal = 16'b0000001011100000;
            15'd5365: log10_cal = 16'b0000001011100000;
            15'd5366: log10_cal = 16'b0000001011100000;
            15'd5367: log10_cal = 16'b0000001011100000;
            15'd5368: log10_cal = 16'b0000001011100000;
            15'd5369: log10_cal = 16'b0000001011100000;
            15'd5370: log10_cal = 16'b0000001011100000;
            15'd5371: log10_cal = 16'b0000001011100001;
            15'd5372: log10_cal = 16'b0000001011100001;
            15'd5373: log10_cal = 16'b0000001011100001;
            15'd5374: log10_cal = 16'b0000001011100001;
            15'd5375: log10_cal = 16'b0000001011100001;
            15'd5376: log10_cal = 16'b0000001011100001;
            15'd5377: log10_cal = 16'b0000001011100001;
            15'd5378: log10_cal = 16'b0000001011100001;
            15'd5379: log10_cal = 16'b0000001011100001;
            15'd5380: log10_cal = 16'b0000001011100001;
            15'd5381: log10_cal = 16'b0000001011100001;
            15'd5382: log10_cal = 16'b0000001011100001;
            15'd5383: log10_cal = 16'b0000001011100010;
            15'd5384: log10_cal = 16'b0000001011100010;
            15'd5385: log10_cal = 16'b0000001011100010;
            15'd5386: log10_cal = 16'b0000001011100010;
            15'd5387: log10_cal = 16'b0000001011100010;
            15'd5388: log10_cal = 16'b0000001011100010;
            15'd5389: log10_cal = 16'b0000001011100010;
            15'd5390: log10_cal = 16'b0000001011100010;
            15'd5391: log10_cal = 16'b0000001011100010;
            15'd5392: log10_cal = 16'b0000001011100010;
            15'd5393: log10_cal = 16'b0000001011100010;
            15'd5394: log10_cal = 16'b0000001011100010;
            15'd5395: log10_cal = 16'b0000001011100011;
            15'd5396: log10_cal = 16'b0000001011100011;
            15'd5397: log10_cal = 16'b0000001011100011;
            15'd5398: log10_cal = 16'b0000001011100011;
            15'd5399: log10_cal = 16'b0000001011100011;
            15'd5400: log10_cal = 16'b0000001011100011;
            15'd5401: log10_cal = 16'b0000001011100011;
            15'd5402: log10_cal = 16'b0000001011100011;
            15'd5403: log10_cal = 16'b0000001011100011;
            15'd5404: log10_cal = 16'b0000001011100011;
            15'd5405: log10_cal = 16'b0000001011100011;
            15'd5406: log10_cal = 16'b0000001011100011;
            15'd5407: log10_cal = 16'b0000001011100100;
            15'd5408: log10_cal = 16'b0000001011100100;
            15'd5409: log10_cal = 16'b0000001011100100;
            15'd5410: log10_cal = 16'b0000001011100100;
            15'd5411: log10_cal = 16'b0000001011100100;
            15'd5412: log10_cal = 16'b0000001011100100;
            15'd5413: log10_cal = 16'b0000001011100100;
            15'd5414: log10_cal = 16'b0000001011100100;
            15'd5415: log10_cal = 16'b0000001011100100;
            15'd5416: log10_cal = 16'b0000001011100100;
            15'd5417: log10_cal = 16'b0000001011100100;
            15'd5418: log10_cal = 16'b0000001011100100;
            15'd5419: log10_cal = 16'b0000001011100100;
            15'd5420: log10_cal = 16'b0000001011100101;
            15'd5421: log10_cal = 16'b0000001011100101;
            15'd5422: log10_cal = 16'b0000001011100101;
            15'd5423: log10_cal = 16'b0000001011100101;
            15'd5424: log10_cal = 16'b0000001011100101;
            15'd5425: log10_cal = 16'b0000001011100101;
            15'd5426: log10_cal = 16'b0000001011100101;
            15'd5427: log10_cal = 16'b0000001011100101;
            15'd5428: log10_cal = 16'b0000001011100101;
            15'd5429: log10_cal = 16'b0000001011100101;
            15'd5430: log10_cal = 16'b0000001011100101;
            15'd5431: log10_cal = 16'b0000001011100101;
            15'd5432: log10_cal = 16'b0000001011100110;
            15'd5433: log10_cal = 16'b0000001011100110;
            15'd5434: log10_cal = 16'b0000001011100110;
            15'd5435: log10_cal = 16'b0000001011100110;
            15'd5436: log10_cal = 16'b0000001011100110;
            15'd5437: log10_cal = 16'b0000001011100110;
            15'd5438: log10_cal = 16'b0000001011100110;
            15'd5439: log10_cal = 16'b0000001011100110;
            15'd5440: log10_cal = 16'b0000001011100110;
            15'd5441: log10_cal = 16'b0000001011100110;
            15'd5442: log10_cal = 16'b0000001011100110;
            15'd5443: log10_cal = 16'b0000001011100110;
            15'd5444: log10_cal = 16'b0000001011100111;
            15'd5445: log10_cal = 16'b0000001011100111;
            15'd5446: log10_cal = 16'b0000001011100111;
            15'd5447: log10_cal = 16'b0000001011100111;
            15'd5448: log10_cal = 16'b0000001011100111;
            15'd5449: log10_cal = 16'b0000001011100111;
            15'd5450: log10_cal = 16'b0000001011100111;
            15'd5451: log10_cal = 16'b0000001011100111;
            15'd5452: log10_cal = 16'b0000001011100111;
            15'd5453: log10_cal = 16'b0000001011100111;
            15'd5454: log10_cal = 16'b0000001011100111;
            15'd5455: log10_cal = 16'b0000001011100111;
            15'd5456: log10_cal = 16'b0000001011101000;
            15'd5457: log10_cal = 16'b0000001011101000;
            15'd5458: log10_cal = 16'b0000001011101000;
            15'd5459: log10_cal = 16'b0000001011101000;
            15'd5460: log10_cal = 16'b0000001011101000;
            15'd5461: log10_cal = 16'b0000001011101000;
            15'd5462: log10_cal = 16'b0000001011101000;
            15'd5463: log10_cal = 16'b0000001011101000;
            15'd5464: log10_cal = 16'b0000001011101000;
            15'd5465: log10_cal = 16'b0000001011101000;
            15'd5466: log10_cal = 16'b0000001011101000;
            15'd5467: log10_cal = 16'b0000001011101000;
            15'd5468: log10_cal = 16'b0000001011101000;
            15'd5469: log10_cal = 16'b0000001011101001;
            15'd5470: log10_cal = 16'b0000001011101001;
            15'd5471: log10_cal = 16'b0000001011101001;
            15'd5472: log10_cal = 16'b0000001011101001;
            15'd5473: log10_cal = 16'b0000001011101001;
            15'd5474: log10_cal = 16'b0000001011101001;
            15'd5475: log10_cal = 16'b0000001011101001;
            15'd5476: log10_cal = 16'b0000001011101001;
            15'd5477: log10_cal = 16'b0000001011101001;
            15'd5478: log10_cal = 16'b0000001011101001;
            15'd5479: log10_cal = 16'b0000001011101001;
            15'd5480: log10_cal = 16'b0000001011101001;
            15'd5481: log10_cal = 16'b0000001011101010;
            15'd5482: log10_cal = 16'b0000001011101010;
            15'd5483: log10_cal = 16'b0000001011101010;
            15'd5484: log10_cal = 16'b0000001011101010;
            15'd5485: log10_cal = 16'b0000001011101010;
            15'd5486: log10_cal = 16'b0000001011101010;
            15'd5487: log10_cal = 16'b0000001011101010;
            15'd5488: log10_cal = 16'b0000001011101010;
            15'd5489: log10_cal = 16'b0000001011101010;
            15'd5490: log10_cal = 16'b0000001011101010;
            15'd5491: log10_cal = 16'b0000001011101010;
            15'd5492: log10_cal = 16'b0000001011101010;
            15'd5493: log10_cal = 16'b0000001011101011;
            15'd5494: log10_cal = 16'b0000001011101011;
            15'd5495: log10_cal = 16'b0000001011101011;
            15'd5496: log10_cal = 16'b0000001011101011;
            15'd5497: log10_cal = 16'b0000001011101011;
            15'd5498: log10_cal = 16'b0000001011101011;
            15'd5499: log10_cal = 16'b0000001011101011;
            15'd5500: log10_cal = 16'b0000001011101011;
            15'd5501: log10_cal = 16'b0000001011101011;
            15'd5502: log10_cal = 16'b0000001011101011;
            15'd5503: log10_cal = 16'b0000001011101011;
            15'd5504: log10_cal = 16'b0000001011101011;
            15'd5505: log10_cal = 16'b0000001011101011;
            15'd5506: log10_cal = 16'b0000001011101100;
            15'd5507: log10_cal = 16'b0000001011101100;
            15'd5508: log10_cal = 16'b0000001011101100;
            15'd5509: log10_cal = 16'b0000001011101100;
            15'd5510: log10_cal = 16'b0000001011101100;
            15'd5511: log10_cal = 16'b0000001011101100;
            15'd5512: log10_cal = 16'b0000001011101100;
            15'd5513: log10_cal = 16'b0000001011101100;
            15'd5514: log10_cal = 16'b0000001011101100;
            15'd5515: log10_cal = 16'b0000001011101100;
            15'd5516: log10_cal = 16'b0000001011101100;
            15'd5517: log10_cal = 16'b0000001011101100;
            15'd5518: log10_cal = 16'b0000001011101101;
            15'd5519: log10_cal = 16'b0000001011101101;
            15'd5520: log10_cal = 16'b0000001011101101;
            15'd5521: log10_cal = 16'b0000001011101101;
            15'd5522: log10_cal = 16'b0000001011101101;
            15'd5523: log10_cal = 16'b0000001011101101;
            15'd5524: log10_cal = 16'b0000001011101101;
            15'd5525: log10_cal = 16'b0000001011101101;
            15'd5526: log10_cal = 16'b0000001011101101;
            15'd5527: log10_cal = 16'b0000001011101101;
            15'd5528: log10_cal = 16'b0000001011101101;
            15'd5529: log10_cal = 16'b0000001011101101;
            15'd5530: log10_cal = 16'b0000001011101110;
            15'd5531: log10_cal = 16'b0000001011101110;
            15'd5532: log10_cal = 16'b0000001011101110;
            15'd5533: log10_cal = 16'b0000001011101110;
            15'd5534: log10_cal = 16'b0000001011101110;
            15'd5535: log10_cal = 16'b0000001011101110;
            15'd5536: log10_cal = 16'b0000001011101110;
            15'd5537: log10_cal = 16'b0000001011101110;
            15'd5538: log10_cal = 16'b0000001011101110;
            15'd5539: log10_cal = 16'b0000001011101110;
            15'd5540: log10_cal = 16'b0000001011101110;
            15'd5541: log10_cal = 16'b0000001011101110;
            15'd5542: log10_cal = 16'b0000001011101110;
            15'd5543: log10_cal = 16'b0000001011101111;
            15'd5544: log10_cal = 16'b0000001011101111;
            15'd5545: log10_cal = 16'b0000001011101111;
            15'd5546: log10_cal = 16'b0000001011101111;
            15'd5547: log10_cal = 16'b0000001011101111;
            15'd5548: log10_cal = 16'b0000001011101111;
            15'd5549: log10_cal = 16'b0000001011101111;
            15'd5550: log10_cal = 16'b0000001011101111;
            15'd5551: log10_cal = 16'b0000001011101111;
            15'd5552: log10_cal = 16'b0000001011101111;
            15'd5553: log10_cal = 16'b0000001011101111;
            15'd5554: log10_cal = 16'b0000001011101111;
            15'd5555: log10_cal = 16'b0000001011110000;
            15'd5556: log10_cal = 16'b0000001011110000;
            15'd5557: log10_cal = 16'b0000001011110000;
            15'd5558: log10_cal = 16'b0000001011110000;
            15'd5559: log10_cal = 16'b0000001011110000;
            15'd5560: log10_cal = 16'b0000001011110000;
            15'd5561: log10_cal = 16'b0000001011110000;
            15'd5562: log10_cal = 16'b0000001011110000;
            15'd5563: log10_cal = 16'b0000001011110000;
            15'd5564: log10_cal = 16'b0000001011110000;
            15'd5565: log10_cal = 16'b0000001011110000;
            15'd5566: log10_cal = 16'b0000001011110000;
            15'd5567: log10_cal = 16'b0000001011110000;
            15'd5568: log10_cal = 16'b0000001011110001;
            15'd5569: log10_cal = 16'b0000001011110001;
            15'd5570: log10_cal = 16'b0000001011110001;
            15'd5571: log10_cal = 16'b0000001011110001;
            15'd5572: log10_cal = 16'b0000001011110001;
            15'd5573: log10_cal = 16'b0000001011110001;
            15'd5574: log10_cal = 16'b0000001011110001;
            15'd5575: log10_cal = 16'b0000001011110001;
            15'd5576: log10_cal = 16'b0000001011110001;
            15'd5577: log10_cal = 16'b0000001011110001;
            15'd5578: log10_cal = 16'b0000001011110001;
            15'd5579: log10_cal = 16'b0000001011110001;
            15'd5580: log10_cal = 16'b0000001011110010;
            15'd5581: log10_cal = 16'b0000001011110010;
            15'd5582: log10_cal = 16'b0000001011110010;
            15'd5583: log10_cal = 16'b0000001011110010;
            15'd5584: log10_cal = 16'b0000001011110010;
            15'd5585: log10_cal = 16'b0000001011110010;
            15'd5586: log10_cal = 16'b0000001011110010;
            15'd5587: log10_cal = 16'b0000001011110010;
            15'd5588: log10_cal = 16'b0000001011110010;
            15'd5589: log10_cal = 16'b0000001011110010;
            15'd5590: log10_cal = 16'b0000001011110010;
            15'd5591: log10_cal = 16'b0000001011110010;
            15'd5592: log10_cal = 16'b0000001011110010;
            15'd5593: log10_cal = 16'b0000001011110011;
            15'd5594: log10_cal = 16'b0000001011110011;
            15'd5595: log10_cal = 16'b0000001011110011;
            15'd5596: log10_cal = 16'b0000001011110011;
            15'd5597: log10_cal = 16'b0000001011110011;
            15'd5598: log10_cal = 16'b0000001011110011;
            15'd5599: log10_cal = 16'b0000001011110011;
            15'd5600: log10_cal = 16'b0000001011110011;
            15'd5601: log10_cal = 16'b0000001011110011;
            15'd5602: log10_cal = 16'b0000001011110011;
            15'd5603: log10_cal = 16'b0000001011110011;
            15'd5604: log10_cal = 16'b0000001011110011;
            15'd5605: log10_cal = 16'b0000001011110011;
            15'd5606: log10_cal = 16'b0000001011110100;
            15'd5607: log10_cal = 16'b0000001011110100;
            15'd5608: log10_cal = 16'b0000001011110100;
            15'd5609: log10_cal = 16'b0000001011110100;
            15'd5610: log10_cal = 16'b0000001011110100;
            15'd5611: log10_cal = 16'b0000001011110100;
            15'd5612: log10_cal = 16'b0000001011110100;
            15'd5613: log10_cal = 16'b0000001011110100;
            15'd5614: log10_cal = 16'b0000001011110100;
            15'd5615: log10_cal = 16'b0000001011110100;
            15'd5616: log10_cal = 16'b0000001011110100;
            15'd5617: log10_cal = 16'b0000001011110100;
            15'd5618: log10_cal = 16'b0000001011110101;
            15'd5619: log10_cal = 16'b0000001011110101;
            15'd5620: log10_cal = 16'b0000001011110101;
            15'd5621: log10_cal = 16'b0000001011110101;
            15'd5622: log10_cal = 16'b0000001011110101;
            15'd5623: log10_cal = 16'b0000001011110101;
            15'd5624: log10_cal = 16'b0000001011110101;
            15'd5625: log10_cal = 16'b0000001011110101;
            15'd5626: log10_cal = 16'b0000001011110101;
            15'd5627: log10_cal = 16'b0000001011110101;
            15'd5628: log10_cal = 16'b0000001011110101;
            15'd5629: log10_cal = 16'b0000001011110101;
            15'd5630: log10_cal = 16'b0000001011110101;
            15'd5631: log10_cal = 16'b0000001011110110;
            15'd5632: log10_cal = 16'b0000001011110110;
            15'd5633: log10_cal = 16'b0000001011110110;
            15'd5634: log10_cal = 16'b0000001011110110;
            15'd5635: log10_cal = 16'b0000001011110110;
            15'd5636: log10_cal = 16'b0000001011110110;
            15'd5637: log10_cal = 16'b0000001011110110;
            15'd5638: log10_cal = 16'b0000001011110110;
            15'd5639: log10_cal = 16'b0000001011110110;
            15'd5640: log10_cal = 16'b0000001011110110;
            15'd5641: log10_cal = 16'b0000001011110110;
            15'd5642: log10_cal = 16'b0000001011110110;
            15'd5643: log10_cal = 16'b0000001011110110;
            15'd5644: log10_cal = 16'b0000001011110111;
            15'd5645: log10_cal = 16'b0000001011110111;
            15'd5646: log10_cal = 16'b0000001011110111;
            15'd5647: log10_cal = 16'b0000001011110111;
            15'd5648: log10_cal = 16'b0000001011110111;
            15'd5649: log10_cal = 16'b0000001011110111;
            15'd5650: log10_cal = 16'b0000001011110111;
            15'd5651: log10_cal = 16'b0000001011110111;
            15'd5652: log10_cal = 16'b0000001011110111;
            15'd5653: log10_cal = 16'b0000001011110111;
            15'd5654: log10_cal = 16'b0000001011110111;
            15'd5655: log10_cal = 16'b0000001011110111;
            15'd5656: log10_cal = 16'b0000001011111000;
            15'd5657: log10_cal = 16'b0000001011111000;
            15'd5658: log10_cal = 16'b0000001011111000;
            15'd5659: log10_cal = 16'b0000001011111000;
            15'd5660: log10_cal = 16'b0000001011111000;
            15'd5661: log10_cal = 16'b0000001011111000;
            15'd5662: log10_cal = 16'b0000001011111000;
            15'd5663: log10_cal = 16'b0000001011111000;
            15'd5664: log10_cal = 16'b0000001011111000;
            15'd5665: log10_cal = 16'b0000001011111000;
            15'd5666: log10_cal = 16'b0000001011111000;
            15'd5667: log10_cal = 16'b0000001011111000;
            15'd5668: log10_cal = 16'b0000001011111000;
            15'd5669: log10_cal = 16'b0000001011111001;
            15'd5670: log10_cal = 16'b0000001011111001;
            15'd5671: log10_cal = 16'b0000001011111001;
            15'd5672: log10_cal = 16'b0000001011111001;
            15'd5673: log10_cal = 16'b0000001011111001;
            15'd5674: log10_cal = 16'b0000001011111001;
            15'd5675: log10_cal = 16'b0000001011111001;
            15'd5676: log10_cal = 16'b0000001011111001;
            15'd5677: log10_cal = 16'b0000001011111001;
            15'd5678: log10_cal = 16'b0000001011111001;
            15'd5679: log10_cal = 16'b0000001011111001;
            15'd5680: log10_cal = 16'b0000001011111001;
            15'd5681: log10_cal = 16'b0000001011111001;
            15'd5682: log10_cal = 16'b0000001011111010;
            15'd5683: log10_cal = 16'b0000001011111010;
            15'd5684: log10_cal = 16'b0000001011111010;
            15'd5685: log10_cal = 16'b0000001011111010;
            15'd5686: log10_cal = 16'b0000001011111010;
            15'd5687: log10_cal = 16'b0000001011111010;
            15'd5688: log10_cal = 16'b0000001011111010;
            15'd5689: log10_cal = 16'b0000001011111010;
            15'd5690: log10_cal = 16'b0000001011111010;
            15'd5691: log10_cal = 16'b0000001011111010;
            15'd5692: log10_cal = 16'b0000001011111010;
            15'd5693: log10_cal = 16'b0000001011111010;
            15'd5694: log10_cal = 16'b0000001011111011;
            15'd5695: log10_cal = 16'b0000001011111011;
            15'd5696: log10_cal = 16'b0000001011111011;
            15'd5697: log10_cal = 16'b0000001011111011;
            15'd5698: log10_cal = 16'b0000001011111011;
            15'd5699: log10_cal = 16'b0000001011111011;
            15'd5700: log10_cal = 16'b0000001011111011;
            15'd5701: log10_cal = 16'b0000001011111011;
            15'd5702: log10_cal = 16'b0000001011111011;
            15'd5703: log10_cal = 16'b0000001011111011;
            15'd5704: log10_cal = 16'b0000001011111011;
            15'd5705: log10_cal = 16'b0000001011111011;
            15'd5706: log10_cal = 16'b0000001011111011;
            15'd5707: log10_cal = 16'b0000001011111100;
            15'd5708: log10_cal = 16'b0000001011111100;
            15'd5709: log10_cal = 16'b0000001011111100;
            15'd5710: log10_cal = 16'b0000001011111100;
            15'd5711: log10_cal = 16'b0000001011111100;
            15'd5712: log10_cal = 16'b0000001011111100;
            15'd5713: log10_cal = 16'b0000001011111100;
            15'd5714: log10_cal = 16'b0000001011111100;
            15'd5715: log10_cal = 16'b0000001011111100;
            15'd5716: log10_cal = 16'b0000001011111100;
            15'd5717: log10_cal = 16'b0000001011111100;
            15'd5718: log10_cal = 16'b0000001011111100;
            15'd5719: log10_cal = 16'b0000001011111100;
            15'd5720: log10_cal = 16'b0000001011111101;
            15'd5721: log10_cal = 16'b0000001011111101;
            15'd5722: log10_cal = 16'b0000001011111101;
            15'd5723: log10_cal = 16'b0000001011111101;
            15'd5724: log10_cal = 16'b0000001011111101;
            15'd5725: log10_cal = 16'b0000001011111101;
            15'd5726: log10_cal = 16'b0000001011111101;
            15'd5727: log10_cal = 16'b0000001011111101;
            15'd5728: log10_cal = 16'b0000001011111101;
            15'd5729: log10_cal = 16'b0000001011111101;
            15'd5730: log10_cal = 16'b0000001011111101;
            15'd5731: log10_cal = 16'b0000001011111101;
            15'd5732: log10_cal = 16'b0000001011111101;
            15'd5733: log10_cal = 16'b0000001011111110;
            15'd5734: log10_cal = 16'b0000001011111110;
            15'd5735: log10_cal = 16'b0000001011111110;
            15'd5736: log10_cal = 16'b0000001011111110;
            15'd5737: log10_cal = 16'b0000001011111110;
            15'd5738: log10_cal = 16'b0000001011111110;
            15'd5739: log10_cal = 16'b0000001011111110;
            15'd5740: log10_cal = 16'b0000001011111110;
            15'd5741: log10_cal = 16'b0000001011111110;
            15'd5742: log10_cal = 16'b0000001011111110;
            15'd5743: log10_cal = 16'b0000001011111110;
            15'd5744: log10_cal = 16'b0000001011111110;
            15'd5745: log10_cal = 16'b0000001011111110;
            15'd5746: log10_cal = 16'b0000001011111111;
            15'd5747: log10_cal = 16'b0000001011111111;
            15'd5748: log10_cal = 16'b0000001011111111;
            15'd5749: log10_cal = 16'b0000001011111111;
            15'd5750: log10_cal = 16'b0000001011111111;
            15'd5751: log10_cal = 16'b0000001011111111;
            15'd5752: log10_cal = 16'b0000001011111111;
            15'd5753: log10_cal = 16'b0000001011111111;
            15'd5754: log10_cal = 16'b0000001011111111;
            15'd5755: log10_cal = 16'b0000001011111111;
            15'd5756: log10_cal = 16'b0000001011111111;
            15'd5757: log10_cal = 16'b0000001011111111;
            15'd5758: log10_cal = 16'b0000001011111111;
            15'd5759: log10_cal = 16'b0000001100000000;
            15'd5760: log10_cal = 16'b0000001100000000;
            15'd5761: log10_cal = 16'b0000001100000000;
            15'd5762: log10_cal = 16'b0000001100000000;
            15'd5763: log10_cal = 16'b0000001100000000;
            15'd5764: log10_cal = 16'b0000001100000000;
            15'd5765: log10_cal = 16'b0000001100000000;
            15'd5766: log10_cal = 16'b0000001100000000;
            15'd5767: log10_cal = 16'b0000001100000000;
            15'd5768: log10_cal = 16'b0000001100000000;
            15'd5769: log10_cal = 16'b0000001100000000;
            15'd5770: log10_cal = 16'b0000001100000000;
            15'd5771: log10_cal = 16'b0000001100000000;
            15'd5772: log10_cal = 16'b0000001100000001;
            15'd5773: log10_cal = 16'b0000001100000001;
            15'd5774: log10_cal = 16'b0000001100000001;
            15'd5775: log10_cal = 16'b0000001100000001;
            15'd5776: log10_cal = 16'b0000001100000001;
            15'd5777: log10_cal = 16'b0000001100000001;
            15'd5778: log10_cal = 16'b0000001100000001;
            15'd5779: log10_cal = 16'b0000001100000001;
            15'd5780: log10_cal = 16'b0000001100000001;
            15'd5781: log10_cal = 16'b0000001100000001;
            15'd5782: log10_cal = 16'b0000001100000001;
            15'd5783: log10_cal = 16'b0000001100000001;
            15'd5784: log10_cal = 16'b0000001100000001;
            15'd5785: log10_cal = 16'b0000001100000010;
            15'd5786: log10_cal = 16'b0000001100000010;
            15'd5787: log10_cal = 16'b0000001100000010;
            15'd5788: log10_cal = 16'b0000001100000010;
            15'd5789: log10_cal = 16'b0000001100000010;
            15'd5790: log10_cal = 16'b0000001100000010;
            15'd5791: log10_cal = 16'b0000001100000010;
            15'd5792: log10_cal = 16'b0000001100000010;
            15'd5793: log10_cal = 16'b0000001100000010;
            15'd5794: log10_cal = 16'b0000001100000010;
            15'd5795: log10_cal = 16'b0000001100000010;
            15'd5796: log10_cal = 16'b0000001100000010;
            15'd5797: log10_cal = 16'b0000001100000010;
            15'd5798: log10_cal = 16'b0000001100000011;
            15'd5799: log10_cal = 16'b0000001100000011;
            15'd5800: log10_cal = 16'b0000001100000011;
            15'd5801: log10_cal = 16'b0000001100000011;
            15'd5802: log10_cal = 16'b0000001100000011;
            15'd5803: log10_cal = 16'b0000001100000011;
            15'd5804: log10_cal = 16'b0000001100000011;
            15'd5805: log10_cal = 16'b0000001100000011;
            15'd5806: log10_cal = 16'b0000001100000011;
            15'd5807: log10_cal = 16'b0000001100000011;
            15'd5808: log10_cal = 16'b0000001100000011;
            15'd5809: log10_cal = 16'b0000001100000011;
            15'd5810: log10_cal = 16'b0000001100000011;
            15'd5811: log10_cal = 16'b0000001100000100;
            15'd5812: log10_cal = 16'b0000001100000100;
            15'd5813: log10_cal = 16'b0000001100000100;
            15'd5814: log10_cal = 16'b0000001100000100;
            15'd5815: log10_cal = 16'b0000001100000100;
            15'd5816: log10_cal = 16'b0000001100000100;
            15'd5817: log10_cal = 16'b0000001100000100;
            15'd5818: log10_cal = 16'b0000001100000100;
            15'd5819: log10_cal = 16'b0000001100000100;
            15'd5820: log10_cal = 16'b0000001100000100;
            15'd5821: log10_cal = 16'b0000001100000100;
            15'd5822: log10_cal = 16'b0000001100000100;
            15'd5823: log10_cal = 16'b0000001100000100;
            15'd5824: log10_cal = 16'b0000001100000101;
            15'd5825: log10_cal = 16'b0000001100000101;
            15'd5826: log10_cal = 16'b0000001100000101;
            15'd5827: log10_cal = 16'b0000001100000101;
            15'd5828: log10_cal = 16'b0000001100000101;
            15'd5829: log10_cal = 16'b0000001100000101;
            15'd5830: log10_cal = 16'b0000001100000101;
            15'd5831: log10_cal = 16'b0000001100000101;
            15'd5832: log10_cal = 16'b0000001100000101;
            15'd5833: log10_cal = 16'b0000001100000101;
            15'd5834: log10_cal = 16'b0000001100000101;
            15'd5835: log10_cal = 16'b0000001100000101;
            15'd5836: log10_cal = 16'b0000001100000101;
            15'd5837: log10_cal = 16'b0000001100000110;
            15'd5838: log10_cal = 16'b0000001100000110;
            15'd5839: log10_cal = 16'b0000001100000110;
            15'd5840: log10_cal = 16'b0000001100000110;
            15'd5841: log10_cal = 16'b0000001100000110;
            15'd5842: log10_cal = 16'b0000001100000110;
            15'd5843: log10_cal = 16'b0000001100000110;
            15'd5844: log10_cal = 16'b0000001100000110;
            15'd5845: log10_cal = 16'b0000001100000110;
            15'd5846: log10_cal = 16'b0000001100000110;
            15'd5847: log10_cal = 16'b0000001100000110;
            15'd5848: log10_cal = 16'b0000001100000110;
            15'd5849: log10_cal = 16'b0000001100000110;
            15'd5850: log10_cal = 16'b0000001100000111;
            15'd5851: log10_cal = 16'b0000001100000111;
            15'd5852: log10_cal = 16'b0000001100000111;
            15'd5853: log10_cal = 16'b0000001100000111;
            15'd5854: log10_cal = 16'b0000001100000111;
            15'd5855: log10_cal = 16'b0000001100000111;
            15'd5856: log10_cal = 16'b0000001100000111;
            15'd5857: log10_cal = 16'b0000001100000111;
            15'd5858: log10_cal = 16'b0000001100000111;
            15'd5859: log10_cal = 16'b0000001100000111;
            15'd5860: log10_cal = 16'b0000001100000111;
            15'd5861: log10_cal = 16'b0000001100000111;
            15'd5862: log10_cal = 16'b0000001100000111;
            15'd5863: log10_cal = 16'b0000001100001000;
            15'd5864: log10_cal = 16'b0000001100001000;
            15'd5865: log10_cal = 16'b0000001100001000;
            15'd5866: log10_cal = 16'b0000001100001000;
            15'd5867: log10_cal = 16'b0000001100001000;
            15'd5868: log10_cal = 16'b0000001100001000;
            15'd5869: log10_cal = 16'b0000001100001000;
            15'd5870: log10_cal = 16'b0000001100001000;
            15'd5871: log10_cal = 16'b0000001100001000;
            15'd5872: log10_cal = 16'b0000001100001000;
            15'd5873: log10_cal = 16'b0000001100001000;
            15'd5874: log10_cal = 16'b0000001100001000;
            15'd5875: log10_cal = 16'b0000001100001000;
            15'd5876: log10_cal = 16'b0000001100001000;
            15'd5877: log10_cal = 16'b0000001100001001;
            15'd5878: log10_cal = 16'b0000001100001001;
            15'd5879: log10_cal = 16'b0000001100001001;
            15'd5880: log10_cal = 16'b0000001100001001;
            15'd5881: log10_cal = 16'b0000001100001001;
            15'd5882: log10_cal = 16'b0000001100001001;
            15'd5883: log10_cal = 16'b0000001100001001;
            15'd5884: log10_cal = 16'b0000001100001001;
            15'd5885: log10_cal = 16'b0000001100001001;
            15'd5886: log10_cal = 16'b0000001100001001;
            15'd5887: log10_cal = 16'b0000001100001001;
            15'd5888: log10_cal = 16'b0000001100001001;
            15'd5889: log10_cal = 16'b0000001100001001;
            15'd5890: log10_cal = 16'b0000001100001010;
            15'd5891: log10_cal = 16'b0000001100001010;
            15'd5892: log10_cal = 16'b0000001100001010;
            15'd5893: log10_cal = 16'b0000001100001010;
            15'd5894: log10_cal = 16'b0000001100001010;
            15'd5895: log10_cal = 16'b0000001100001010;
            15'd5896: log10_cal = 16'b0000001100001010;
            15'd5897: log10_cal = 16'b0000001100001010;
            15'd5898: log10_cal = 16'b0000001100001010;
            15'd5899: log10_cal = 16'b0000001100001010;
            15'd5900: log10_cal = 16'b0000001100001010;
            15'd5901: log10_cal = 16'b0000001100001010;
            15'd5902: log10_cal = 16'b0000001100001010;
            15'd5903: log10_cal = 16'b0000001100001011;
            15'd5904: log10_cal = 16'b0000001100001011;
            15'd5905: log10_cal = 16'b0000001100001011;
            15'd5906: log10_cal = 16'b0000001100001011;
            15'd5907: log10_cal = 16'b0000001100001011;
            15'd5908: log10_cal = 16'b0000001100001011;
            15'd5909: log10_cal = 16'b0000001100001011;
            15'd5910: log10_cal = 16'b0000001100001011;
            15'd5911: log10_cal = 16'b0000001100001011;
            15'd5912: log10_cal = 16'b0000001100001011;
            15'd5913: log10_cal = 16'b0000001100001011;
            15'd5914: log10_cal = 16'b0000001100001011;
            15'd5915: log10_cal = 16'b0000001100001011;
            15'd5916: log10_cal = 16'b0000001100001100;
            15'd5917: log10_cal = 16'b0000001100001100;
            15'd5918: log10_cal = 16'b0000001100001100;
            15'd5919: log10_cal = 16'b0000001100001100;
            15'd5920: log10_cal = 16'b0000001100001100;
            15'd5921: log10_cal = 16'b0000001100001100;
            15'd5922: log10_cal = 16'b0000001100001100;
            15'd5923: log10_cal = 16'b0000001100001100;
            15'd5924: log10_cal = 16'b0000001100001100;
            15'd5925: log10_cal = 16'b0000001100001100;
            15'd5926: log10_cal = 16'b0000001100001100;
            15'd5927: log10_cal = 16'b0000001100001100;
            15'd5928: log10_cal = 16'b0000001100001100;
            15'd5929: log10_cal = 16'b0000001100001100;
            15'd5930: log10_cal = 16'b0000001100001101;
            15'd5931: log10_cal = 16'b0000001100001101;
            15'd5932: log10_cal = 16'b0000001100001101;
            15'd5933: log10_cal = 16'b0000001100001101;
            15'd5934: log10_cal = 16'b0000001100001101;
            15'd5935: log10_cal = 16'b0000001100001101;
            15'd5936: log10_cal = 16'b0000001100001101;
            15'd5937: log10_cal = 16'b0000001100001101;
            15'd5938: log10_cal = 16'b0000001100001101;
            15'd5939: log10_cal = 16'b0000001100001101;
            15'd5940: log10_cal = 16'b0000001100001101;
            15'd5941: log10_cal = 16'b0000001100001101;
            15'd5942: log10_cal = 16'b0000001100001101;
            15'd5943: log10_cal = 16'b0000001100001110;
            15'd5944: log10_cal = 16'b0000001100001110;
            15'd5945: log10_cal = 16'b0000001100001110;
            15'd5946: log10_cal = 16'b0000001100001110;
            15'd5947: log10_cal = 16'b0000001100001110;
            15'd5948: log10_cal = 16'b0000001100001110;
            15'd5949: log10_cal = 16'b0000001100001110;
            15'd5950: log10_cal = 16'b0000001100001110;
            15'd5951: log10_cal = 16'b0000001100001110;
            15'd5952: log10_cal = 16'b0000001100001110;
            15'd5953: log10_cal = 16'b0000001100001110;
            15'd5954: log10_cal = 16'b0000001100001110;
            15'd5955: log10_cal = 16'b0000001100001110;
            15'd5956: log10_cal = 16'b0000001100001111;
            15'd5957: log10_cal = 16'b0000001100001111;
            15'd5958: log10_cal = 16'b0000001100001111;
            15'd5959: log10_cal = 16'b0000001100001111;
            15'd5960: log10_cal = 16'b0000001100001111;
            15'd5961: log10_cal = 16'b0000001100001111;
            15'd5962: log10_cal = 16'b0000001100001111;
            15'd5963: log10_cal = 16'b0000001100001111;
            15'd5964: log10_cal = 16'b0000001100001111;
            15'd5965: log10_cal = 16'b0000001100001111;
            15'd5966: log10_cal = 16'b0000001100001111;
            15'd5967: log10_cal = 16'b0000001100001111;
            15'd5968: log10_cal = 16'b0000001100001111;
            15'd5969: log10_cal = 16'b0000001100001111;
            15'd5970: log10_cal = 16'b0000001100010000;
            15'd5971: log10_cal = 16'b0000001100010000;
            15'd5972: log10_cal = 16'b0000001100010000;
            15'd5973: log10_cal = 16'b0000001100010000;
            15'd5974: log10_cal = 16'b0000001100010000;
            15'd5975: log10_cal = 16'b0000001100010000;
            15'd5976: log10_cal = 16'b0000001100010000;
            15'd5977: log10_cal = 16'b0000001100010000;
            15'd5978: log10_cal = 16'b0000001100010000;
            15'd5979: log10_cal = 16'b0000001100010000;
            15'd5980: log10_cal = 16'b0000001100010000;
            15'd5981: log10_cal = 16'b0000001100010000;
            15'd5982: log10_cal = 16'b0000001100010000;
            15'd5983: log10_cal = 16'b0000001100010001;
            15'd5984: log10_cal = 16'b0000001100010001;
            15'd5985: log10_cal = 16'b0000001100010001;
            15'd5986: log10_cal = 16'b0000001100010001;
            15'd5987: log10_cal = 16'b0000001100010001;
            15'd5988: log10_cal = 16'b0000001100010001;
            15'd5989: log10_cal = 16'b0000001100010001;
            15'd5990: log10_cal = 16'b0000001100010001;
            15'd5991: log10_cal = 16'b0000001100010001;
            15'd5992: log10_cal = 16'b0000001100010001;
            15'd5993: log10_cal = 16'b0000001100010001;
            15'd5994: log10_cal = 16'b0000001100010001;
            15'd5995: log10_cal = 16'b0000001100010001;
            15'd5996: log10_cal = 16'b0000001100010001;
            15'd5997: log10_cal = 16'b0000001100010010;
            15'd5998: log10_cal = 16'b0000001100010010;
            15'd5999: log10_cal = 16'b0000001100010010;
            15'd6000: log10_cal = 16'b0000001100010010;
            15'd6001: log10_cal = 16'b0000001100010010;
            15'd6002: log10_cal = 16'b0000001100010010;
            15'd6003: log10_cal = 16'b0000001100010010;
            15'd6004: log10_cal = 16'b0000001100010010;
            15'd6005: log10_cal = 16'b0000001100010010;
            15'd6006: log10_cal = 16'b0000001100010010;
            15'd6007: log10_cal = 16'b0000001100010010;
            15'd6008: log10_cal = 16'b0000001100010010;
            15'd6009: log10_cal = 16'b0000001100010010;
            15'd6010: log10_cal = 16'b0000001100010011;
            15'd6011: log10_cal = 16'b0000001100010011;
            15'd6012: log10_cal = 16'b0000001100010011;
            15'd6013: log10_cal = 16'b0000001100010011;
            15'd6014: log10_cal = 16'b0000001100010011;
            15'd6015: log10_cal = 16'b0000001100010011;
            15'd6016: log10_cal = 16'b0000001100010011;
            15'd6017: log10_cal = 16'b0000001100010011;
            15'd6018: log10_cal = 16'b0000001100010011;
            15'd6019: log10_cal = 16'b0000001100010011;
            15'd6020: log10_cal = 16'b0000001100010011;
            15'd6021: log10_cal = 16'b0000001100010011;
            15'd6022: log10_cal = 16'b0000001100010011;
            15'd6023: log10_cal = 16'b0000001100010011;
            15'd6024: log10_cal = 16'b0000001100010100;
            15'd6025: log10_cal = 16'b0000001100010100;
            15'd6026: log10_cal = 16'b0000001100010100;
            15'd6027: log10_cal = 16'b0000001100010100;
            15'd6028: log10_cal = 16'b0000001100010100;
            15'd6029: log10_cal = 16'b0000001100010100;
            15'd6030: log10_cal = 16'b0000001100010100;
            15'd6031: log10_cal = 16'b0000001100010100;
            15'd6032: log10_cal = 16'b0000001100010100;
            15'd6033: log10_cal = 16'b0000001100010100;
            15'd6034: log10_cal = 16'b0000001100010100;
            15'd6035: log10_cal = 16'b0000001100010100;
            15'd6036: log10_cal = 16'b0000001100010100;
            15'd6037: log10_cal = 16'b0000001100010101;
            15'd6038: log10_cal = 16'b0000001100010101;
            15'd6039: log10_cal = 16'b0000001100010101;
            15'd6040: log10_cal = 16'b0000001100010101;
            15'd6041: log10_cal = 16'b0000001100010101;
            15'd6042: log10_cal = 16'b0000001100010101;
            15'd6043: log10_cal = 16'b0000001100010101;
            15'd6044: log10_cal = 16'b0000001100010101;
            15'd6045: log10_cal = 16'b0000001100010101;
            15'd6046: log10_cal = 16'b0000001100010101;
            15'd6047: log10_cal = 16'b0000001100010101;
            15'd6048: log10_cal = 16'b0000001100010101;
            15'd6049: log10_cal = 16'b0000001100010101;
            15'd6050: log10_cal = 16'b0000001100010101;
            15'd6051: log10_cal = 16'b0000001100010110;
            15'd6052: log10_cal = 16'b0000001100010110;
            15'd6053: log10_cal = 16'b0000001100010110;
            15'd6054: log10_cal = 16'b0000001100010110;
            15'd6055: log10_cal = 16'b0000001100010110;
            15'd6056: log10_cal = 16'b0000001100010110;
            15'd6057: log10_cal = 16'b0000001100010110;
            15'd6058: log10_cal = 16'b0000001100010110;
            15'd6059: log10_cal = 16'b0000001100010110;
            15'd6060: log10_cal = 16'b0000001100010110;
            15'd6061: log10_cal = 16'b0000001100010110;
            15'd6062: log10_cal = 16'b0000001100010110;
            15'd6063: log10_cal = 16'b0000001100010110;
            15'd6064: log10_cal = 16'b0000001100010110;
            15'd6065: log10_cal = 16'b0000001100010111;
            15'd6066: log10_cal = 16'b0000001100010111;
            15'd6067: log10_cal = 16'b0000001100010111;
            15'd6068: log10_cal = 16'b0000001100010111;
            15'd6069: log10_cal = 16'b0000001100010111;
            15'd6070: log10_cal = 16'b0000001100010111;
            15'd6071: log10_cal = 16'b0000001100010111;
            15'd6072: log10_cal = 16'b0000001100010111;
            15'd6073: log10_cal = 16'b0000001100010111;
            15'd6074: log10_cal = 16'b0000001100010111;
            15'd6075: log10_cal = 16'b0000001100010111;
            15'd6076: log10_cal = 16'b0000001100010111;
            15'd6077: log10_cal = 16'b0000001100010111;
            15'd6078: log10_cal = 16'b0000001100011000;
            15'd6079: log10_cal = 16'b0000001100011000;
            15'd6080: log10_cal = 16'b0000001100011000;
            15'd6081: log10_cal = 16'b0000001100011000;
            15'd6082: log10_cal = 16'b0000001100011000;
            15'd6083: log10_cal = 16'b0000001100011000;
            15'd6084: log10_cal = 16'b0000001100011000;
            15'd6085: log10_cal = 16'b0000001100011000;
            15'd6086: log10_cal = 16'b0000001100011000;
            15'd6087: log10_cal = 16'b0000001100011000;
            15'd6088: log10_cal = 16'b0000001100011000;
            15'd6089: log10_cal = 16'b0000001100011000;
            15'd6090: log10_cal = 16'b0000001100011000;
            15'd6091: log10_cal = 16'b0000001100011000;
            15'd6092: log10_cal = 16'b0000001100011001;
            15'd6093: log10_cal = 16'b0000001100011001;
            15'd6094: log10_cal = 16'b0000001100011001;
            15'd6095: log10_cal = 16'b0000001100011001;
            15'd6096: log10_cal = 16'b0000001100011001;
            15'd6097: log10_cal = 16'b0000001100011001;
            15'd6098: log10_cal = 16'b0000001100011001;
            15'd6099: log10_cal = 16'b0000001100011001;
            15'd6100: log10_cal = 16'b0000001100011001;
            15'd6101: log10_cal = 16'b0000001100011001;
            15'd6102: log10_cal = 16'b0000001100011001;
            15'd6103: log10_cal = 16'b0000001100011001;
            15'd6104: log10_cal = 16'b0000001100011001;
            15'd6105: log10_cal = 16'b0000001100011001;
            15'd6106: log10_cal = 16'b0000001100011010;
            15'd6107: log10_cal = 16'b0000001100011010;
            15'd6108: log10_cal = 16'b0000001100011010;
            15'd6109: log10_cal = 16'b0000001100011010;
            15'd6110: log10_cal = 16'b0000001100011010;
            15'd6111: log10_cal = 16'b0000001100011010;
            15'd6112: log10_cal = 16'b0000001100011010;
            15'd6113: log10_cal = 16'b0000001100011010;
            15'd6114: log10_cal = 16'b0000001100011010;
            15'd6115: log10_cal = 16'b0000001100011010;
            15'd6116: log10_cal = 16'b0000001100011010;
            15'd6117: log10_cal = 16'b0000001100011010;
            15'd6118: log10_cal = 16'b0000001100011010;
            15'd6119: log10_cal = 16'b0000001100011011;
            15'd6120: log10_cal = 16'b0000001100011011;
            15'd6121: log10_cal = 16'b0000001100011011;
            15'd6122: log10_cal = 16'b0000001100011011;
            15'd6123: log10_cal = 16'b0000001100011011;
            15'd6124: log10_cal = 16'b0000001100011011;
            15'd6125: log10_cal = 16'b0000001100011011;
            15'd6126: log10_cal = 16'b0000001100011011;
            15'd6127: log10_cal = 16'b0000001100011011;
            15'd6128: log10_cal = 16'b0000001100011011;
            15'd6129: log10_cal = 16'b0000001100011011;
            15'd6130: log10_cal = 16'b0000001100011011;
            15'd6131: log10_cal = 16'b0000001100011011;
            15'd6132: log10_cal = 16'b0000001100011011;
            15'd6133: log10_cal = 16'b0000001100011100;
            15'd6134: log10_cal = 16'b0000001100011100;
            15'd6135: log10_cal = 16'b0000001100011100;
            15'd6136: log10_cal = 16'b0000001100011100;
            15'd6137: log10_cal = 16'b0000001100011100;
            15'd6138: log10_cal = 16'b0000001100011100;
            15'd6139: log10_cal = 16'b0000001100011100;
            15'd6140: log10_cal = 16'b0000001100011100;
            15'd6141: log10_cal = 16'b0000001100011100;
            15'd6142: log10_cal = 16'b0000001100011100;
            15'd6143: log10_cal = 16'b0000001100011100;
            15'd6144: log10_cal = 16'b0000001100011100;
            15'd6145: log10_cal = 16'b0000001100011100;
            15'd6146: log10_cal = 16'b0000001100011100;
            15'd6147: log10_cal = 16'b0000001100011101;
            15'd6148: log10_cal = 16'b0000001100011101;
            15'd6149: log10_cal = 16'b0000001100011101;
            15'd6150: log10_cal = 16'b0000001100011101;
            15'd6151: log10_cal = 16'b0000001100011101;
            15'd6152: log10_cal = 16'b0000001100011101;
            15'd6153: log10_cal = 16'b0000001100011101;
            15'd6154: log10_cal = 16'b0000001100011101;
            15'd6155: log10_cal = 16'b0000001100011101;
            15'd6156: log10_cal = 16'b0000001100011101;
            15'd6157: log10_cal = 16'b0000001100011101;
            15'd6158: log10_cal = 16'b0000001100011101;
            15'd6159: log10_cal = 16'b0000001100011101;
            15'd6160: log10_cal = 16'b0000001100011101;
            15'd6161: log10_cal = 16'b0000001100011110;
            15'd6162: log10_cal = 16'b0000001100011110;
            15'd6163: log10_cal = 16'b0000001100011110;
            15'd6164: log10_cal = 16'b0000001100011110;
            15'd6165: log10_cal = 16'b0000001100011110;
            15'd6166: log10_cal = 16'b0000001100011110;
            15'd6167: log10_cal = 16'b0000001100011110;
            15'd6168: log10_cal = 16'b0000001100011110;
            15'd6169: log10_cal = 16'b0000001100011110;
            15'd6170: log10_cal = 16'b0000001100011110;
            15'd6171: log10_cal = 16'b0000001100011110;
            15'd6172: log10_cal = 16'b0000001100011110;
            15'd6173: log10_cal = 16'b0000001100011110;
            15'd6174: log10_cal = 16'b0000001100011110;
            15'd6175: log10_cal = 16'b0000001100011111;
            15'd6176: log10_cal = 16'b0000001100011111;
            15'd6177: log10_cal = 16'b0000001100011111;
            15'd6178: log10_cal = 16'b0000001100011111;
            15'd6179: log10_cal = 16'b0000001100011111;
            15'd6180: log10_cal = 16'b0000001100011111;
            15'd6181: log10_cal = 16'b0000001100011111;
            15'd6182: log10_cal = 16'b0000001100011111;
            15'd6183: log10_cal = 16'b0000001100011111;
            15'd6184: log10_cal = 16'b0000001100011111;
            15'd6185: log10_cal = 16'b0000001100011111;
            15'd6186: log10_cal = 16'b0000001100011111;
            15'd6187: log10_cal = 16'b0000001100011111;
            15'd6188: log10_cal = 16'b0000001100100000;
            15'd6189: log10_cal = 16'b0000001100100000;
            15'd6190: log10_cal = 16'b0000001100100000;
            15'd6191: log10_cal = 16'b0000001100100000;
            15'd6192: log10_cal = 16'b0000001100100000;
            15'd6193: log10_cal = 16'b0000001100100000;
            15'd6194: log10_cal = 16'b0000001100100000;
            15'd6195: log10_cal = 16'b0000001100100000;
            15'd6196: log10_cal = 16'b0000001100100000;
            15'd6197: log10_cal = 16'b0000001100100000;
            15'd6198: log10_cal = 16'b0000001100100000;
            15'd6199: log10_cal = 16'b0000001100100000;
            15'd6200: log10_cal = 16'b0000001100100000;
            15'd6201: log10_cal = 16'b0000001100100000;
            15'd6202: log10_cal = 16'b0000001100100001;
            15'd6203: log10_cal = 16'b0000001100100001;
            15'd6204: log10_cal = 16'b0000001100100001;
            15'd6205: log10_cal = 16'b0000001100100001;
            15'd6206: log10_cal = 16'b0000001100100001;
            15'd6207: log10_cal = 16'b0000001100100001;
            15'd6208: log10_cal = 16'b0000001100100001;
            15'd6209: log10_cal = 16'b0000001100100001;
            15'd6210: log10_cal = 16'b0000001100100001;
            15'd6211: log10_cal = 16'b0000001100100001;
            15'd6212: log10_cal = 16'b0000001100100001;
            15'd6213: log10_cal = 16'b0000001100100001;
            15'd6214: log10_cal = 16'b0000001100100001;
            15'd6215: log10_cal = 16'b0000001100100001;
            15'd6216: log10_cal = 16'b0000001100100010;
            15'd6217: log10_cal = 16'b0000001100100010;
            15'd6218: log10_cal = 16'b0000001100100010;
            15'd6219: log10_cal = 16'b0000001100100010;
            15'd6220: log10_cal = 16'b0000001100100010;
            15'd6221: log10_cal = 16'b0000001100100010;
            15'd6222: log10_cal = 16'b0000001100100010;
            15'd6223: log10_cal = 16'b0000001100100010;
            15'd6224: log10_cal = 16'b0000001100100010;
            15'd6225: log10_cal = 16'b0000001100100010;
            15'd6226: log10_cal = 16'b0000001100100010;
            15'd6227: log10_cal = 16'b0000001100100010;
            15'd6228: log10_cal = 16'b0000001100100010;
            15'd6229: log10_cal = 16'b0000001100100010;
            15'd6230: log10_cal = 16'b0000001100100011;
            15'd6231: log10_cal = 16'b0000001100100011;
            15'd6232: log10_cal = 16'b0000001100100011;
            15'd6233: log10_cal = 16'b0000001100100011;
            15'd6234: log10_cal = 16'b0000001100100011;
            15'd6235: log10_cal = 16'b0000001100100011;
            15'd6236: log10_cal = 16'b0000001100100011;
            15'd6237: log10_cal = 16'b0000001100100011;
            15'd6238: log10_cal = 16'b0000001100100011;
            15'd6239: log10_cal = 16'b0000001100100011;
            15'd6240: log10_cal = 16'b0000001100100011;
            15'd6241: log10_cal = 16'b0000001100100011;
            15'd6242: log10_cal = 16'b0000001100100011;
            15'd6243: log10_cal = 16'b0000001100100011;
            15'd6244: log10_cal = 16'b0000001100100100;
            15'd6245: log10_cal = 16'b0000001100100100;
            15'd6246: log10_cal = 16'b0000001100100100;
            15'd6247: log10_cal = 16'b0000001100100100;
            15'd6248: log10_cal = 16'b0000001100100100;
            15'd6249: log10_cal = 16'b0000001100100100;
            15'd6250: log10_cal = 16'b0000001100100100;
            15'd6251: log10_cal = 16'b0000001100100100;
            15'd6252: log10_cal = 16'b0000001100100100;
            15'd6253: log10_cal = 16'b0000001100100100;
            15'd6254: log10_cal = 16'b0000001100100100;
            15'd6255: log10_cal = 16'b0000001100100100;
            15'd6256: log10_cal = 16'b0000001100100100;
            15'd6257: log10_cal = 16'b0000001100100100;
            15'd6258: log10_cal = 16'b0000001100100101;
            15'd6259: log10_cal = 16'b0000001100100101;
            15'd6260: log10_cal = 16'b0000001100100101;
            15'd6261: log10_cal = 16'b0000001100100101;
            15'd6262: log10_cal = 16'b0000001100100101;
            15'd6263: log10_cal = 16'b0000001100100101;
            15'd6264: log10_cal = 16'b0000001100100101;
            15'd6265: log10_cal = 16'b0000001100100101;
            15'd6266: log10_cal = 16'b0000001100100101;
            15'd6267: log10_cal = 16'b0000001100100101;
            15'd6268: log10_cal = 16'b0000001100100101;
            15'd6269: log10_cal = 16'b0000001100100101;
            15'd6270: log10_cal = 16'b0000001100100101;
            15'd6271: log10_cal = 16'b0000001100100101;
            15'd6272: log10_cal = 16'b0000001100100101;
            15'd6273: log10_cal = 16'b0000001100100110;
            15'd6274: log10_cal = 16'b0000001100100110;
            15'd6275: log10_cal = 16'b0000001100100110;
            15'd6276: log10_cal = 16'b0000001100100110;
            15'd6277: log10_cal = 16'b0000001100100110;
            15'd6278: log10_cal = 16'b0000001100100110;
            15'd6279: log10_cal = 16'b0000001100100110;
            15'd6280: log10_cal = 16'b0000001100100110;
            15'd6281: log10_cal = 16'b0000001100100110;
            15'd6282: log10_cal = 16'b0000001100100110;
            15'd6283: log10_cal = 16'b0000001100100110;
            15'd6284: log10_cal = 16'b0000001100100110;
            15'd6285: log10_cal = 16'b0000001100100110;
            15'd6286: log10_cal = 16'b0000001100100110;
            15'd6287: log10_cal = 16'b0000001100100111;
            15'd6288: log10_cal = 16'b0000001100100111;
            15'd6289: log10_cal = 16'b0000001100100111;
            15'd6290: log10_cal = 16'b0000001100100111;
            15'd6291: log10_cal = 16'b0000001100100111;
            15'd6292: log10_cal = 16'b0000001100100111;
            15'd6293: log10_cal = 16'b0000001100100111;
            15'd6294: log10_cal = 16'b0000001100100111;
            15'd6295: log10_cal = 16'b0000001100100111;
            15'd6296: log10_cal = 16'b0000001100100111;
            15'd6297: log10_cal = 16'b0000001100100111;
            15'd6298: log10_cal = 16'b0000001100100111;
            15'd6299: log10_cal = 16'b0000001100100111;
            15'd6300: log10_cal = 16'b0000001100100111;
            15'd6301: log10_cal = 16'b0000001100101000;
            15'd6302: log10_cal = 16'b0000001100101000;
            15'd6303: log10_cal = 16'b0000001100101000;
            15'd6304: log10_cal = 16'b0000001100101000;
            15'd6305: log10_cal = 16'b0000001100101000;
            15'd6306: log10_cal = 16'b0000001100101000;
            15'd6307: log10_cal = 16'b0000001100101000;
            15'd6308: log10_cal = 16'b0000001100101000;
            15'd6309: log10_cal = 16'b0000001100101000;
            15'd6310: log10_cal = 16'b0000001100101000;
            15'd6311: log10_cal = 16'b0000001100101000;
            15'd6312: log10_cal = 16'b0000001100101000;
            15'd6313: log10_cal = 16'b0000001100101000;
            15'd6314: log10_cal = 16'b0000001100101000;
            15'd6315: log10_cal = 16'b0000001100101001;
            15'd6316: log10_cal = 16'b0000001100101001;
            15'd6317: log10_cal = 16'b0000001100101001;
            15'd6318: log10_cal = 16'b0000001100101001;
            15'd6319: log10_cal = 16'b0000001100101001;
            15'd6320: log10_cal = 16'b0000001100101001;
            15'd6321: log10_cal = 16'b0000001100101001;
            15'd6322: log10_cal = 16'b0000001100101001;
            15'd6323: log10_cal = 16'b0000001100101001;
            15'd6324: log10_cal = 16'b0000001100101001;
            15'd6325: log10_cal = 16'b0000001100101001;
            15'd6326: log10_cal = 16'b0000001100101001;
            15'd6327: log10_cal = 16'b0000001100101001;
            15'd6328: log10_cal = 16'b0000001100101001;
            15'd6329: log10_cal = 16'b0000001100101010;
            15'd6330: log10_cal = 16'b0000001100101010;
            15'd6331: log10_cal = 16'b0000001100101010;
            15'd6332: log10_cal = 16'b0000001100101010;
            15'd6333: log10_cal = 16'b0000001100101010;
            15'd6334: log10_cal = 16'b0000001100101010;
            15'd6335: log10_cal = 16'b0000001100101010;
            15'd6336: log10_cal = 16'b0000001100101010;
            15'd6337: log10_cal = 16'b0000001100101010;
            15'd6338: log10_cal = 16'b0000001100101010;
            15'd6339: log10_cal = 16'b0000001100101010;
            15'd6340: log10_cal = 16'b0000001100101010;
            15'd6341: log10_cal = 16'b0000001100101010;
            15'd6342: log10_cal = 16'b0000001100101010;
            15'd6343: log10_cal = 16'b0000001100101011;
            15'd6344: log10_cal = 16'b0000001100101011;
            15'd6345: log10_cal = 16'b0000001100101011;
            15'd6346: log10_cal = 16'b0000001100101011;
            15'd6347: log10_cal = 16'b0000001100101011;
            15'd6348: log10_cal = 16'b0000001100101011;
            15'd6349: log10_cal = 16'b0000001100101011;
            15'd6350: log10_cal = 16'b0000001100101011;
            15'd6351: log10_cal = 16'b0000001100101011;
            15'd6352: log10_cal = 16'b0000001100101011;
            15'd6353: log10_cal = 16'b0000001100101011;
            15'd6354: log10_cal = 16'b0000001100101011;
            15'd6355: log10_cal = 16'b0000001100101011;
            15'd6356: log10_cal = 16'b0000001100101011;
            15'd6357: log10_cal = 16'b0000001100101011;
            15'd6358: log10_cal = 16'b0000001100101100;
            15'd6359: log10_cal = 16'b0000001100101100;
            15'd6360: log10_cal = 16'b0000001100101100;
            15'd6361: log10_cal = 16'b0000001100101100;
            15'd6362: log10_cal = 16'b0000001100101100;
            15'd6363: log10_cal = 16'b0000001100101100;
            15'd6364: log10_cal = 16'b0000001100101100;
            15'd6365: log10_cal = 16'b0000001100101100;
            15'd6366: log10_cal = 16'b0000001100101100;
            15'd6367: log10_cal = 16'b0000001100101100;
            15'd6368: log10_cal = 16'b0000001100101100;
            15'd6369: log10_cal = 16'b0000001100101100;
            15'd6370: log10_cal = 16'b0000001100101100;
            15'd6371: log10_cal = 16'b0000001100101100;
            15'd6372: log10_cal = 16'b0000001100101101;
            15'd6373: log10_cal = 16'b0000001100101101;
            15'd6374: log10_cal = 16'b0000001100101101;
            15'd6375: log10_cal = 16'b0000001100101101;
            15'd6376: log10_cal = 16'b0000001100101101;
            15'd6377: log10_cal = 16'b0000001100101101;
            15'd6378: log10_cal = 16'b0000001100101101;
            15'd6379: log10_cal = 16'b0000001100101101;
            15'd6380: log10_cal = 16'b0000001100101101;
            15'd6381: log10_cal = 16'b0000001100101101;
            15'd6382: log10_cal = 16'b0000001100101101;
            15'd6383: log10_cal = 16'b0000001100101101;
            15'd6384: log10_cal = 16'b0000001100101101;
            15'd6385: log10_cal = 16'b0000001100101101;
            15'd6386: log10_cal = 16'b0000001100101110;
            15'd6387: log10_cal = 16'b0000001100101110;
            15'd6388: log10_cal = 16'b0000001100101110;
            15'd6389: log10_cal = 16'b0000001100101110;
            15'd6390: log10_cal = 16'b0000001100101110;
            15'd6391: log10_cal = 16'b0000001100101110;
            15'd6392: log10_cal = 16'b0000001100101110;
            15'd6393: log10_cal = 16'b0000001100101110;
            15'd6394: log10_cal = 16'b0000001100101110;
            15'd6395: log10_cal = 16'b0000001100101110;
            15'd6396: log10_cal = 16'b0000001100101110;
            15'd6397: log10_cal = 16'b0000001100101110;
            15'd6398: log10_cal = 16'b0000001100101110;
            15'd6399: log10_cal = 16'b0000001100101110;
            15'd6400: log10_cal = 16'b0000001100101110;
            15'd6401: log10_cal = 16'b0000001100101111;
            15'd6402: log10_cal = 16'b0000001100101111;
            15'd6403: log10_cal = 16'b0000001100101111;
            15'd6404: log10_cal = 16'b0000001100101111;
            15'd6405: log10_cal = 16'b0000001100101111;
            15'd6406: log10_cal = 16'b0000001100101111;
            15'd6407: log10_cal = 16'b0000001100101111;
            15'd6408: log10_cal = 16'b0000001100101111;
            15'd6409: log10_cal = 16'b0000001100101111;
            15'd6410: log10_cal = 16'b0000001100101111;
            15'd6411: log10_cal = 16'b0000001100101111;
            15'd6412: log10_cal = 16'b0000001100101111;
            15'd6413: log10_cal = 16'b0000001100101111;
            15'd6414: log10_cal = 16'b0000001100101111;
            15'd6415: log10_cal = 16'b0000001100110000;
            15'd6416: log10_cal = 16'b0000001100110000;
            15'd6417: log10_cal = 16'b0000001100110000;
            15'd6418: log10_cal = 16'b0000001100110000;
            15'd6419: log10_cal = 16'b0000001100110000;
            15'd6420: log10_cal = 16'b0000001100110000;
            15'd6421: log10_cal = 16'b0000001100110000;
            15'd6422: log10_cal = 16'b0000001100110000;
            15'd6423: log10_cal = 16'b0000001100110000;
            15'd6424: log10_cal = 16'b0000001100110000;
            15'd6425: log10_cal = 16'b0000001100110000;
            15'd6426: log10_cal = 16'b0000001100110000;
            15'd6427: log10_cal = 16'b0000001100110000;
            15'd6428: log10_cal = 16'b0000001100110000;
            15'd6429: log10_cal = 16'b0000001100110000;
            15'd6430: log10_cal = 16'b0000001100110001;
            15'd6431: log10_cal = 16'b0000001100110001;
            15'd6432: log10_cal = 16'b0000001100110001;
            15'd6433: log10_cal = 16'b0000001100110001;
            15'd6434: log10_cal = 16'b0000001100110001;
            15'd6435: log10_cal = 16'b0000001100110001;
            15'd6436: log10_cal = 16'b0000001100110001;
            15'd6437: log10_cal = 16'b0000001100110001;
            15'd6438: log10_cal = 16'b0000001100110001;
            15'd6439: log10_cal = 16'b0000001100110001;
            15'd6440: log10_cal = 16'b0000001100110001;
            15'd6441: log10_cal = 16'b0000001100110001;
            15'd6442: log10_cal = 16'b0000001100110001;
            15'd6443: log10_cal = 16'b0000001100110001;
            15'd6444: log10_cal = 16'b0000001100110010;
            15'd6445: log10_cal = 16'b0000001100110010;
            15'd6446: log10_cal = 16'b0000001100110010;
            15'd6447: log10_cal = 16'b0000001100110010;
            15'd6448: log10_cal = 16'b0000001100110010;
            15'd6449: log10_cal = 16'b0000001100110010;
            15'd6450: log10_cal = 16'b0000001100110010;
            15'd6451: log10_cal = 16'b0000001100110010;
            15'd6452: log10_cal = 16'b0000001100110010;
            15'd6453: log10_cal = 16'b0000001100110010;
            15'd6454: log10_cal = 16'b0000001100110010;
            15'd6455: log10_cal = 16'b0000001100110010;
            15'd6456: log10_cal = 16'b0000001100110010;
            15'd6457: log10_cal = 16'b0000001100110010;
            15'd6458: log10_cal = 16'b0000001100110010;
            15'd6459: log10_cal = 16'b0000001100110011;
            15'd6460: log10_cal = 16'b0000001100110011;
            15'd6461: log10_cal = 16'b0000001100110011;
            15'd6462: log10_cal = 16'b0000001100110011;
            15'd6463: log10_cal = 16'b0000001100110011;
            15'd6464: log10_cal = 16'b0000001100110011;
            15'd6465: log10_cal = 16'b0000001100110011;
            15'd6466: log10_cal = 16'b0000001100110011;
            15'd6467: log10_cal = 16'b0000001100110011;
            15'd6468: log10_cal = 16'b0000001100110011;
            15'd6469: log10_cal = 16'b0000001100110011;
            15'd6470: log10_cal = 16'b0000001100110011;
            15'd6471: log10_cal = 16'b0000001100110011;
            15'd6472: log10_cal = 16'b0000001100110011;
            15'd6473: log10_cal = 16'b0000001100110100;
            15'd6474: log10_cal = 16'b0000001100110100;
            15'd6475: log10_cal = 16'b0000001100110100;
            15'd6476: log10_cal = 16'b0000001100110100;
            15'd6477: log10_cal = 16'b0000001100110100;
            15'd6478: log10_cal = 16'b0000001100110100;
            15'd6479: log10_cal = 16'b0000001100110100;
            15'd6480: log10_cal = 16'b0000001100110100;
            15'd6481: log10_cal = 16'b0000001100110100;
            15'd6482: log10_cal = 16'b0000001100110100;
            15'd6483: log10_cal = 16'b0000001100110100;
            15'd6484: log10_cal = 16'b0000001100110100;
            15'd6485: log10_cal = 16'b0000001100110100;
            15'd6486: log10_cal = 16'b0000001100110100;
            15'd6487: log10_cal = 16'b0000001100110100;
            15'd6488: log10_cal = 16'b0000001100110101;
            15'd6489: log10_cal = 16'b0000001100110101;
            15'd6490: log10_cal = 16'b0000001100110101;
            15'd6491: log10_cal = 16'b0000001100110101;
            15'd6492: log10_cal = 16'b0000001100110101;
            15'd6493: log10_cal = 16'b0000001100110101;
            15'd6494: log10_cal = 16'b0000001100110101;
            15'd6495: log10_cal = 16'b0000001100110101;
            15'd6496: log10_cal = 16'b0000001100110101;
            15'd6497: log10_cal = 16'b0000001100110101;
            15'd6498: log10_cal = 16'b0000001100110101;
            15'd6499: log10_cal = 16'b0000001100110101;
            15'd6500: log10_cal = 16'b0000001100110101;
            15'd6501: log10_cal = 16'b0000001100110101;
            15'd6502: log10_cal = 16'b0000001100110110;
            15'd6503: log10_cal = 16'b0000001100110110;
            15'd6504: log10_cal = 16'b0000001100110110;
            15'd6505: log10_cal = 16'b0000001100110110;
            15'd6506: log10_cal = 16'b0000001100110110;
            15'd6507: log10_cal = 16'b0000001100110110;
            15'd6508: log10_cal = 16'b0000001100110110;
            15'd6509: log10_cal = 16'b0000001100110110;
            15'd6510: log10_cal = 16'b0000001100110110;
            15'd6511: log10_cal = 16'b0000001100110110;
            15'd6512: log10_cal = 16'b0000001100110110;
            15'd6513: log10_cal = 16'b0000001100110110;
            15'd6514: log10_cal = 16'b0000001100110110;
            15'd6515: log10_cal = 16'b0000001100110110;
            15'd6516: log10_cal = 16'b0000001100110110;
            15'd6517: log10_cal = 16'b0000001100110111;
            15'd6518: log10_cal = 16'b0000001100110111;
            15'd6519: log10_cal = 16'b0000001100110111;
            15'd6520: log10_cal = 16'b0000001100110111;
            15'd6521: log10_cal = 16'b0000001100110111;
            15'd6522: log10_cal = 16'b0000001100110111;
            15'd6523: log10_cal = 16'b0000001100110111;
            15'd6524: log10_cal = 16'b0000001100110111;
            15'd6525: log10_cal = 16'b0000001100110111;
            15'd6526: log10_cal = 16'b0000001100110111;
            15'd6527: log10_cal = 16'b0000001100110111;
            15'd6528: log10_cal = 16'b0000001100110111;
            15'd6529: log10_cal = 16'b0000001100110111;
            15'd6530: log10_cal = 16'b0000001100110111;
            15'd6531: log10_cal = 16'b0000001100110111;
            15'd6532: log10_cal = 16'b0000001100111000;
            15'd6533: log10_cal = 16'b0000001100111000;
            15'd6534: log10_cal = 16'b0000001100111000;
            15'd6535: log10_cal = 16'b0000001100111000;
            15'd6536: log10_cal = 16'b0000001100111000;
            15'd6537: log10_cal = 16'b0000001100111000;
            15'd6538: log10_cal = 16'b0000001100111000;
            15'd6539: log10_cal = 16'b0000001100111000;
            15'd6540: log10_cal = 16'b0000001100111000;
            15'd6541: log10_cal = 16'b0000001100111000;
            15'd6542: log10_cal = 16'b0000001100111000;
            15'd6543: log10_cal = 16'b0000001100111000;
            15'd6544: log10_cal = 16'b0000001100111000;
            15'd6545: log10_cal = 16'b0000001100111000;
            15'd6546: log10_cal = 16'b0000001100111001;
            15'd6547: log10_cal = 16'b0000001100111001;
            15'd6548: log10_cal = 16'b0000001100111001;
            15'd6549: log10_cal = 16'b0000001100111001;
            15'd6550: log10_cal = 16'b0000001100111001;
            15'd6551: log10_cal = 16'b0000001100111001;
            15'd6552: log10_cal = 16'b0000001100111001;
            15'd6553: log10_cal = 16'b0000001100111001;
            15'd6554: log10_cal = 16'b0000001100111001;
            15'd6555: log10_cal = 16'b0000001100111001;
            15'd6556: log10_cal = 16'b0000001100111001;
            15'd6557: log10_cal = 16'b0000001100111001;
            15'd6558: log10_cal = 16'b0000001100111001;
            15'd6559: log10_cal = 16'b0000001100111001;
            15'd6560: log10_cal = 16'b0000001100111001;
            15'd6561: log10_cal = 16'b0000001100111010;
            15'd6562: log10_cal = 16'b0000001100111010;
            15'd6563: log10_cal = 16'b0000001100111010;
            15'd6564: log10_cal = 16'b0000001100111010;
            15'd6565: log10_cal = 16'b0000001100111010;
            15'd6566: log10_cal = 16'b0000001100111010;
            15'd6567: log10_cal = 16'b0000001100111010;
            15'd6568: log10_cal = 16'b0000001100111010;
            15'd6569: log10_cal = 16'b0000001100111010;
            15'd6570: log10_cal = 16'b0000001100111010;
            15'd6571: log10_cal = 16'b0000001100111010;
            15'd6572: log10_cal = 16'b0000001100111010;
            15'd6573: log10_cal = 16'b0000001100111010;
            15'd6574: log10_cal = 16'b0000001100111010;
            15'd6575: log10_cal = 16'b0000001100111010;
            15'd6576: log10_cal = 16'b0000001100111011;
            15'd6577: log10_cal = 16'b0000001100111011;
            15'd6578: log10_cal = 16'b0000001100111011;
            15'd6579: log10_cal = 16'b0000001100111011;
            15'd6580: log10_cal = 16'b0000001100111011;
            15'd6581: log10_cal = 16'b0000001100111011;
            15'd6582: log10_cal = 16'b0000001100111011;
            15'd6583: log10_cal = 16'b0000001100111011;
            15'd6584: log10_cal = 16'b0000001100111011;
            15'd6585: log10_cal = 16'b0000001100111011;
            15'd6586: log10_cal = 16'b0000001100111011;
            15'd6587: log10_cal = 16'b0000001100111011;
            15'd6588: log10_cal = 16'b0000001100111011;
            15'd6589: log10_cal = 16'b0000001100111011;
            15'd6590: log10_cal = 16'b0000001100111011;
            15'd6591: log10_cal = 16'b0000001100111100;
            15'd6592: log10_cal = 16'b0000001100111100;
            15'd6593: log10_cal = 16'b0000001100111100;
            15'd6594: log10_cal = 16'b0000001100111100;
            15'd6595: log10_cal = 16'b0000001100111100;
            15'd6596: log10_cal = 16'b0000001100111100;
            15'd6597: log10_cal = 16'b0000001100111100;
            15'd6598: log10_cal = 16'b0000001100111100;
            15'd6599: log10_cal = 16'b0000001100111100;
            15'd6600: log10_cal = 16'b0000001100111100;
            15'd6601: log10_cal = 16'b0000001100111100;
            15'd6602: log10_cal = 16'b0000001100111100;
            15'd6603: log10_cal = 16'b0000001100111100;
            15'd6604: log10_cal = 16'b0000001100111100;
            15'd6605: log10_cal = 16'b0000001100111101;
            15'd6606: log10_cal = 16'b0000001100111101;
            15'd6607: log10_cal = 16'b0000001100111101;
            15'd6608: log10_cal = 16'b0000001100111101;
            15'd6609: log10_cal = 16'b0000001100111101;
            15'd6610: log10_cal = 16'b0000001100111101;
            15'd6611: log10_cal = 16'b0000001100111101;
            15'd6612: log10_cal = 16'b0000001100111101;
            15'd6613: log10_cal = 16'b0000001100111101;
            15'd6614: log10_cal = 16'b0000001100111101;
            15'd6615: log10_cal = 16'b0000001100111101;
            15'd6616: log10_cal = 16'b0000001100111101;
            15'd6617: log10_cal = 16'b0000001100111101;
            15'd6618: log10_cal = 16'b0000001100111101;
            15'd6619: log10_cal = 16'b0000001100111101;
            15'd6620: log10_cal = 16'b0000001100111110;
            15'd6621: log10_cal = 16'b0000001100111110;
            15'd6622: log10_cal = 16'b0000001100111110;
            15'd6623: log10_cal = 16'b0000001100111110;
            15'd6624: log10_cal = 16'b0000001100111110;
            15'd6625: log10_cal = 16'b0000001100111110;
            15'd6626: log10_cal = 16'b0000001100111110;
            15'd6627: log10_cal = 16'b0000001100111110;
            15'd6628: log10_cal = 16'b0000001100111110;
            15'd6629: log10_cal = 16'b0000001100111110;
            15'd6630: log10_cal = 16'b0000001100111110;
            15'd6631: log10_cal = 16'b0000001100111110;
            15'd6632: log10_cal = 16'b0000001100111110;
            15'd6633: log10_cal = 16'b0000001100111110;
            15'd6634: log10_cal = 16'b0000001100111110;
            15'd6635: log10_cal = 16'b0000001100111111;
            15'd6636: log10_cal = 16'b0000001100111111;
            15'd6637: log10_cal = 16'b0000001100111111;
            15'd6638: log10_cal = 16'b0000001100111111;
            15'd6639: log10_cal = 16'b0000001100111111;
            15'd6640: log10_cal = 16'b0000001100111111;
            15'd6641: log10_cal = 16'b0000001100111111;
            15'd6642: log10_cal = 16'b0000001100111111;
            15'd6643: log10_cal = 16'b0000001100111111;
            15'd6644: log10_cal = 16'b0000001100111111;
            15'd6645: log10_cal = 16'b0000001100111111;
            15'd6646: log10_cal = 16'b0000001100111111;
            15'd6647: log10_cal = 16'b0000001100111111;
            15'd6648: log10_cal = 16'b0000001100111111;
            15'd6649: log10_cal = 16'b0000001100111111;
            15'd6650: log10_cal = 16'b0000001101000000;
            15'd6651: log10_cal = 16'b0000001101000000;
            15'd6652: log10_cal = 16'b0000001101000000;
            15'd6653: log10_cal = 16'b0000001101000000;
            15'd6654: log10_cal = 16'b0000001101000000;
            15'd6655: log10_cal = 16'b0000001101000000;
            15'd6656: log10_cal = 16'b0000001101000000;
            15'd6657: log10_cal = 16'b0000001101000000;
            15'd6658: log10_cal = 16'b0000001101000000;
            15'd6659: log10_cal = 16'b0000001101000000;
            15'd6660: log10_cal = 16'b0000001101000000;
            15'd6661: log10_cal = 16'b0000001101000000;
            15'd6662: log10_cal = 16'b0000001101000000;
            15'd6663: log10_cal = 16'b0000001101000000;
            15'd6664: log10_cal = 16'b0000001101000000;
            15'd6665: log10_cal = 16'b0000001101000001;
            15'd6666: log10_cal = 16'b0000001101000001;
            15'd6667: log10_cal = 16'b0000001101000001;
            15'd6668: log10_cal = 16'b0000001101000001;
            15'd6669: log10_cal = 16'b0000001101000001;
            15'd6670: log10_cal = 16'b0000001101000001;
            15'd6671: log10_cal = 16'b0000001101000001;
            15'd6672: log10_cal = 16'b0000001101000001;
            15'd6673: log10_cal = 16'b0000001101000001;
            15'd6674: log10_cal = 16'b0000001101000001;
            15'd6675: log10_cal = 16'b0000001101000001;
            15'd6676: log10_cal = 16'b0000001101000001;
            15'd6677: log10_cal = 16'b0000001101000001;
            15'd6678: log10_cal = 16'b0000001101000001;
            15'd6679: log10_cal = 16'b0000001101000001;
            15'd6680: log10_cal = 16'b0000001101000010;
            15'd6681: log10_cal = 16'b0000001101000010;
            15'd6682: log10_cal = 16'b0000001101000010;
            15'd6683: log10_cal = 16'b0000001101000010;
            15'd6684: log10_cal = 16'b0000001101000010;
            15'd6685: log10_cal = 16'b0000001101000010;
            15'd6686: log10_cal = 16'b0000001101000010;
            15'd6687: log10_cal = 16'b0000001101000010;
            15'd6688: log10_cal = 16'b0000001101000010;
            15'd6689: log10_cal = 16'b0000001101000010;
            15'd6690: log10_cal = 16'b0000001101000010;
            15'd6691: log10_cal = 16'b0000001101000010;
            15'd6692: log10_cal = 16'b0000001101000010;
            15'd6693: log10_cal = 16'b0000001101000010;
            15'd6694: log10_cal = 16'b0000001101000010;
            15'd6695: log10_cal = 16'b0000001101000011;
            15'd6696: log10_cal = 16'b0000001101000011;
            15'd6697: log10_cal = 16'b0000001101000011;
            15'd6698: log10_cal = 16'b0000001101000011;
            15'd6699: log10_cal = 16'b0000001101000011;
            15'd6700: log10_cal = 16'b0000001101000011;
            15'd6701: log10_cal = 16'b0000001101000011;
            15'd6702: log10_cal = 16'b0000001101000011;
            15'd6703: log10_cal = 16'b0000001101000011;
            15'd6704: log10_cal = 16'b0000001101000011;
            15'd6705: log10_cal = 16'b0000001101000011;
            15'd6706: log10_cal = 16'b0000001101000011;
            15'd6707: log10_cal = 16'b0000001101000011;
            15'd6708: log10_cal = 16'b0000001101000011;
            15'd6709: log10_cal = 16'b0000001101000011;
            15'd6710: log10_cal = 16'b0000001101000100;
            15'd6711: log10_cal = 16'b0000001101000100;
            15'd6712: log10_cal = 16'b0000001101000100;
            15'd6713: log10_cal = 16'b0000001101000100;
            15'd6714: log10_cal = 16'b0000001101000100;
            15'd6715: log10_cal = 16'b0000001101000100;
            15'd6716: log10_cal = 16'b0000001101000100;
            15'd6717: log10_cal = 16'b0000001101000100;
            15'd6718: log10_cal = 16'b0000001101000100;
            15'd6719: log10_cal = 16'b0000001101000100;
            15'd6720: log10_cal = 16'b0000001101000100;
            15'd6721: log10_cal = 16'b0000001101000100;
            15'd6722: log10_cal = 16'b0000001101000100;
            15'd6723: log10_cal = 16'b0000001101000100;
            15'd6724: log10_cal = 16'b0000001101000100;
            15'd6725: log10_cal = 16'b0000001101000101;
            15'd6726: log10_cal = 16'b0000001101000101;
            15'd6727: log10_cal = 16'b0000001101000101;
            15'd6728: log10_cal = 16'b0000001101000101;
            15'd6729: log10_cal = 16'b0000001101000101;
            15'd6730: log10_cal = 16'b0000001101000101;
            15'd6731: log10_cal = 16'b0000001101000101;
            15'd6732: log10_cal = 16'b0000001101000101;
            15'd6733: log10_cal = 16'b0000001101000101;
            15'd6734: log10_cal = 16'b0000001101000101;
            15'd6735: log10_cal = 16'b0000001101000101;
            15'd6736: log10_cal = 16'b0000001101000101;
            15'd6737: log10_cal = 16'b0000001101000101;
            15'd6738: log10_cal = 16'b0000001101000101;
            15'd6739: log10_cal = 16'b0000001101000101;
            15'd6740: log10_cal = 16'b0000001101000110;
            15'd6741: log10_cal = 16'b0000001101000110;
            15'd6742: log10_cal = 16'b0000001101000110;
            15'd6743: log10_cal = 16'b0000001101000110;
            15'd6744: log10_cal = 16'b0000001101000110;
            15'd6745: log10_cal = 16'b0000001101000110;
            15'd6746: log10_cal = 16'b0000001101000110;
            15'd6747: log10_cal = 16'b0000001101000110;
            15'd6748: log10_cal = 16'b0000001101000110;
            15'd6749: log10_cal = 16'b0000001101000110;
            15'd6750: log10_cal = 16'b0000001101000110;
            15'd6751: log10_cal = 16'b0000001101000110;
            15'd6752: log10_cal = 16'b0000001101000110;
            15'd6753: log10_cal = 16'b0000001101000110;
            15'd6754: log10_cal = 16'b0000001101000110;
            15'd6755: log10_cal = 16'b0000001101000110;
            15'd6756: log10_cal = 16'b0000001101000111;
            15'd6757: log10_cal = 16'b0000001101000111;
            15'd6758: log10_cal = 16'b0000001101000111;
            15'd6759: log10_cal = 16'b0000001101000111;
            15'd6760: log10_cal = 16'b0000001101000111;
            15'd6761: log10_cal = 16'b0000001101000111;
            15'd6762: log10_cal = 16'b0000001101000111;
            15'd6763: log10_cal = 16'b0000001101000111;
            15'd6764: log10_cal = 16'b0000001101000111;
            15'd6765: log10_cal = 16'b0000001101000111;
            15'd6766: log10_cal = 16'b0000001101000111;
            15'd6767: log10_cal = 16'b0000001101000111;
            15'd6768: log10_cal = 16'b0000001101000111;
            15'd6769: log10_cal = 16'b0000001101000111;
            15'd6770: log10_cal = 16'b0000001101000111;
            15'd6771: log10_cal = 16'b0000001101001000;
            15'd6772: log10_cal = 16'b0000001101001000;
            15'd6773: log10_cal = 16'b0000001101001000;
            15'd6774: log10_cal = 16'b0000001101001000;
            15'd6775: log10_cal = 16'b0000001101001000;
            15'd6776: log10_cal = 16'b0000001101001000;
            15'd6777: log10_cal = 16'b0000001101001000;
            15'd6778: log10_cal = 16'b0000001101001000;
            15'd6779: log10_cal = 16'b0000001101001000;
            15'd6780: log10_cal = 16'b0000001101001000;
            15'd6781: log10_cal = 16'b0000001101001000;
            15'd6782: log10_cal = 16'b0000001101001000;
            15'd6783: log10_cal = 16'b0000001101001000;
            15'd6784: log10_cal = 16'b0000001101001000;
            15'd6785: log10_cal = 16'b0000001101001000;
            15'd6786: log10_cal = 16'b0000001101001001;
            15'd6787: log10_cal = 16'b0000001101001001;
            15'd6788: log10_cal = 16'b0000001101001001;
            15'd6789: log10_cal = 16'b0000001101001001;
            15'd6790: log10_cal = 16'b0000001101001001;
            15'd6791: log10_cal = 16'b0000001101001001;
            15'd6792: log10_cal = 16'b0000001101001001;
            15'd6793: log10_cal = 16'b0000001101001001;
            15'd6794: log10_cal = 16'b0000001101001001;
            15'd6795: log10_cal = 16'b0000001101001001;
            15'd6796: log10_cal = 16'b0000001101001001;
            15'd6797: log10_cal = 16'b0000001101001001;
            15'd6798: log10_cal = 16'b0000001101001001;
            15'd6799: log10_cal = 16'b0000001101001001;
            15'd6800: log10_cal = 16'b0000001101001001;
            15'd6801: log10_cal = 16'b0000001101001010;
            15'd6802: log10_cal = 16'b0000001101001010;
            15'd6803: log10_cal = 16'b0000001101001010;
            15'd6804: log10_cal = 16'b0000001101001010;
            15'd6805: log10_cal = 16'b0000001101001010;
            15'd6806: log10_cal = 16'b0000001101001010;
            15'd6807: log10_cal = 16'b0000001101001010;
            15'd6808: log10_cal = 16'b0000001101001010;
            15'd6809: log10_cal = 16'b0000001101001010;
            15'd6810: log10_cal = 16'b0000001101001010;
            15'd6811: log10_cal = 16'b0000001101001010;
            15'd6812: log10_cal = 16'b0000001101001010;
            15'd6813: log10_cal = 16'b0000001101001010;
            15'd6814: log10_cal = 16'b0000001101001010;
            15'd6815: log10_cal = 16'b0000001101001010;
            15'd6816: log10_cal = 16'b0000001101001010;
            15'd6817: log10_cal = 16'b0000001101001011;
            15'd6818: log10_cal = 16'b0000001101001011;
            15'd6819: log10_cal = 16'b0000001101001011;
            15'd6820: log10_cal = 16'b0000001101001011;
            15'd6821: log10_cal = 16'b0000001101001011;
            15'd6822: log10_cal = 16'b0000001101001011;
            15'd6823: log10_cal = 16'b0000001101001011;
            15'd6824: log10_cal = 16'b0000001101001011;
            15'd6825: log10_cal = 16'b0000001101001011;
            15'd6826: log10_cal = 16'b0000001101001011;
            15'd6827: log10_cal = 16'b0000001101001011;
            15'd6828: log10_cal = 16'b0000001101001011;
            15'd6829: log10_cal = 16'b0000001101001011;
            15'd6830: log10_cal = 16'b0000001101001011;
            15'd6831: log10_cal = 16'b0000001101001011;
            15'd6832: log10_cal = 16'b0000001101001100;
            15'd6833: log10_cal = 16'b0000001101001100;
            15'd6834: log10_cal = 16'b0000001101001100;
            15'd6835: log10_cal = 16'b0000001101001100;
            15'd6836: log10_cal = 16'b0000001101001100;
            15'd6837: log10_cal = 16'b0000001101001100;
            15'd6838: log10_cal = 16'b0000001101001100;
            15'd6839: log10_cal = 16'b0000001101001100;
            15'd6840: log10_cal = 16'b0000001101001100;
            15'd6841: log10_cal = 16'b0000001101001100;
            15'd6842: log10_cal = 16'b0000001101001100;
            15'd6843: log10_cal = 16'b0000001101001100;
            15'd6844: log10_cal = 16'b0000001101001100;
            15'd6845: log10_cal = 16'b0000001101001100;
            15'd6846: log10_cal = 16'b0000001101001100;
            15'd6847: log10_cal = 16'b0000001101001101;
            15'd6848: log10_cal = 16'b0000001101001101;
            15'd6849: log10_cal = 16'b0000001101001101;
            15'd6850: log10_cal = 16'b0000001101001101;
            15'd6851: log10_cal = 16'b0000001101001101;
            15'd6852: log10_cal = 16'b0000001101001101;
            15'd6853: log10_cal = 16'b0000001101001101;
            15'd6854: log10_cal = 16'b0000001101001101;
            15'd6855: log10_cal = 16'b0000001101001101;
            15'd6856: log10_cal = 16'b0000001101001101;
            15'd6857: log10_cal = 16'b0000001101001101;
            15'd6858: log10_cal = 16'b0000001101001101;
            15'd6859: log10_cal = 16'b0000001101001101;
            15'd6860: log10_cal = 16'b0000001101001101;
            15'd6861: log10_cal = 16'b0000001101001101;
            15'd6862: log10_cal = 16'b0000001101001101;
            15'd6863: log10_cal = 16'b0000001101001110;
            15'd6864: log10_cal = 16'b0000001101001110;
            15'd6865: log10_cal = 16'b0000001101001110;
            15'd6866: log10_cal = 16'b0000001101001110;
            15'd6867: log10_cal = 16'b0000001101001110;
            15'd6868: log10_cal = 16'b0000001101001110;
            15'd6869: log10_cal = 16'b0000001101001110;
            15'd6870: log10_cal = 16'b0000001101001110;
            15'd6871: log10_cal = 16'b0000001101001110;
            15'd6872: log10_cal = 16'b0000001101001110;
            15'd6873: log10_cal = 16'b0000001101001110;
            15'd6874: log10_cal = 16'b0000001101001110;
            15'd6875: log10_cal = 16'b0000001101001110;
            15'd6876: log10_cal = 16'b0000001101001110;
            15'd6877: log10_cal = 16'b0000001101001110;
            15'd6878: log10_cal = 16'b0000001101001111;
            15'd6879: log10_cal = 16'b0000001101001111;
            15'd6880: log10_cal = 16'b0000001101001111;
            15'd6881: log10_cal = 16'b0000001101001111;
            15'd6882: log10_cal = 16'b0000001101001111;
            15'd6883: log10_cal = 16'b0000001101001111;
            15'd6884: log10_cal = 16'b0000001101001111;
            15'd6885: log10_cal = 16'b0000001101001111;
            15'd6886: log10_cal = 16'b0000001101001111;
            15'd6887: log10_cal = 16'b0000001101001111;
            15'd6888: log10_cal = 16'b0000001101001111;
            15'd6889: log10_cal = 16'b0000001101001111;
            15'd6890: log10_cal = 16'b0000001101001111;
            15'd6891: log10_cal = 16'b0000001101001111;
            15'd6892: log10_cal = 16'b0000001101001111;
            15'd6893: log10_cal = 16'b0000001101001111;
            15'd6894: log10_cal = 16'b0000001101010000;
            15'd6895: log10_cal = 16'b0000001101010000;
            15'd6896: log10_cal = 16'b0000001101010000;
            15'd6897: log10_cal = 16'b0000001101010000;
            15'd6898: log10_cal = 16'b0000001101010000;
            15'd6899: log10_cal = 16'b0000001101010000;
            15'd6900: log10_cal = 16'b0000001101010000;
            15'd6901: log10_cal = 16'b0000001101010000;
            15'd6902: log10_cal = 16'b0000001101010000;
            15'd6903: log10_cal = 16'b0000001101010000;
            15'd6904: log10_cal = 16'b0000001101010000;
            15'd6905: log10_cal = 16'b0000001101010000;
            15'd6906: log10_cal = 16'b0000001101010000;
            15'd6907: log10_cal = 16'b0000001101010000;
            15'd6908: log10_cal = 16'b0000001101010000;
            15'd6909: log10_cal = 16'b0000001101010001;
            15'd6910: log10_cal = 16'b0000001101010001;
            15'd6911: log10_cal = 16'b0000001101010001;
            15'd6912: log10_cal = 16'b0000001101010001;
            15'd6913: log10_cal = 16'b0000001101010001;
            15'd6914: log10_cal = 16'b0000001101010001;
            15'd6915: log10_cal = 16'b0000001101010001;
            15'd6916: log10_cal = 16'b0000001101010001;
            15'd6917: log10_cal = 16'b0000001101010001;
            15'd6918: log10_cal = 16'b0000001101010001;
            15'd6919: log10_cal = 16'b0000001101010001;
            15'd6920: log10_cal = 16'b0000001101010001;
            15'd6921: log10_cal = 16'b0000001101010001;
            15'd6922: log10_cal = 16'b0000001101010001;
            15'd6923: log10_cal = 16'b0000001101010001;
            15'd6924: log10_cal = 16'b0000001101010001;
            15'd6925: log10_cal = 16'b0000001101010010;
            15'd6926: log10_cal = 16'b0000001101010010;
            15'd6927: log10_cal = 16'b0000001101010010;
            15'd6928: log10_cal = 16'b0000001101010010;
            15'd6929: log10_cal = 16'b0000001101010010;
            15'd6930: log10_cal = 16'b0000001101010010;
            15'd6931: log10_cal = 16'b0000001101010010;
            15'd6932: log10_cal = 16'b0000001101010010;
            15'd6933: log10_cal = 16'b0000001101010010;
            15'd6934: log10_cal = 16'b0000001101010010;
            15'd6935: log10_cal = 16'b0000001101010010;
            15'd6936: log10_cal = 16'b0000001101010010;
            15'd6937: log10_cal = 16'b0000001101010010;
            15'd6938: log10_cal = 16'b0000001101010010;
            15'd6939: log10_cal = 16'b0000001101010010;
            15'd6940: log10_cal = 16'b0000001101010011;
            15'd6941: log10_cal = 16'b0000001101010011;
            15'd6942: log10_cal = 16'b0000001101010011;
            15'd6943: log10_cal = 16'b0000001101010011;
            15'd6944: log10_cal = 16'b0000001101010011;
            15'd6945: log10_cal = 16'b0000001101010011;
            15'd6946: log10_cal = 16'b0000001101010011;
            15'd6947: log10_cal = 16'b0000001101010011;
            15'd6948: log10_cal = 16'b0000001101010011;
            15'd6949: log10_cal = 16'b0000001101010011;
            15'd6950: log10_cal = 16'b0000001101010011;
            15'd6951: log10_cal = 16'b0000001101010011;
            15'd6952: log10_cal = 16'b0000001101010011;
            15'd6953: log10_cal = 16'b0000001101010011;
            15'd6954: log10_cal = 16'b0000001101010011;
            15'd6955: log10_cal = 16'b0000001101010011;
            15'd6956: log10_cal = 16'b0000001101010100;
            15'd6957: log10_cal = 16'b0000001101010100;
            15'd6958: log10_cal = 16'b0000001101010100;
            15'd6959: log10_cal = 16'b0000001101010100;
            15'd6960: log10_cal = 16'b0000001101010100;
            15'd6961: log10_cal = 16'b0000001101010100;
            15'd6962: log10_cal = 16'b0000001101010100;
            15'd6963: log10_cal = 16'b0000001101010100;
            15'd6964: log10_cal = 16'b0000001101010100;
            15'd6965: log10_cal = 16'b0000001101010100;
            15'd6966: log10_cal = 16'b0000001101010100;
            15'd6967: log10_cal = 16'b0000001101010100;
            15'd6968: log10_cal = 16'b0000001101010100;
            15'd6969: log10_cal = 16'b0000001101010100;
            15'd6970: log10_cal = 16'b0000001101010100;
            15'd6971: log10_cal = 16'b0000001101010100;
            15'd6972: log10_cal = 16'b0000001101010101;
            15'd6973: log10_cal = 16'b0000001101010101;
            15'd6974: log10_cal = 16'b0000001101010101;
            15'd6975: log10_cal = 16'b0000001101010101;
            15'd6976: log10_cal = 16'b0000001101010101;
            15'd6977: log10_cal = 16'b0000001101010101;
            15'd6978: log10_cal = 16'b0000001101010101;
            15'd6979: log10_cal = 16'b0000001101010101;
            15'd6980: log10_cal = 16'b0000001101010101;
            15'd6981: log10_cal = 16'b0000001101010101;
            15'd6982: log10_cal = 16'b0000001101010101;
            15'd6983: log10_cal = 16'b0000001101010101;
            15'd6984: log10_cal = 16'b0000001101010101;
            15'd6985: log10_cal = 16'b0000001101010101;
            15'd6986: log10_cal = 16'b0000001101010101;
            15'd6987: log10_cal = 16'b0000001101010110;
            15'd6988: log10_cal = 16'b0000001101010110;
            15'd6989: log10_cal = 16'b0000001101010110;
            15'd6990: log10_cal = 16'b0000001101010110;
            15'd6991: log10_cal = 16'b0000001101010110;
            15'd6992: log10_cal = 16'b0000001101010110;
            15'd6993: log10_cal = 16'b0000001101010110;
            15'd6994: log10_cal = 16'b0000001101010110;
            15'd6995: log10_cal = 16'b0000001101010110;
            15'd6996: log10_cal = 16'b0000001101010110;
            15'd6997: log10_cal = 16'b0000001101010110;
            15'd6998: log10_cal = 16'b0000001101010110;
            15'd6999: log10_cal = 16'b0000001101010110;
            15'd7000: log10_cal = 16'b0000001101010110;
            15'd7001: log10_cal = 16'b0000001101010110;
            15'd7002: log10_cal = 16'b0000001101010110;
            15'd7003: log10_cal = 16'b0000001101010111;
            15'd7004: log10_cal = 16'b0000001101010111;
            15'd7005: log10_cal = 16'b0000001101010111;
            15'd7006: log10_cal = 16'b0000001101010111;
            15'd7007: log10_cal = 16'b0000001101010111;
            15'd7008: log10_cal = 16'b0000001101010111;
            15'd7009: log10_cal = 16'b0000001101010111;
            15'd7010: log10_cal = 16'b0000001101010111;
            15'd7011: log10_cal = 16'b0000001101010111;
            15'd7012: log10_cal = 16'b0000001101010111;
            15'd7013: log10_cal = 16'b0000001101010111;
            15'd7014: log10_cal = 16'b0000001101010111;
            15'd7015: log10_cal = 16'b0000001101010111;
            15'd7016: log10_cal = 16'b0000001101010111;
            15'd7017: log10_cal = 16'b0000001101010111;
            15'd7018: log10_cal = 16'b0000001101010111;
            15'd7019: log10_cal = 16'b0000001101011000;
            15'd7020: log10_cal = 16'b0000001101011000;
            15'd7021: log10_cal = 16'b0000001101011000;
            15'd7022: log10_cal = 16'b0000001101011000;
            15'd7023: log10_cal = 16'b0000001101011000;
            15'd7024: log10_cal = 16'b0000001101011000;
            15'd7025: log10_cal = 16'b0000001101011000;
            15'd7026: log10_cal = 16'b0000001101011000;
            15'd7027: log10_cal = 16'b0000001101011000;
            15'd7028: log10_cal = 16'b0000001101011000;
            15'd7029: log10_cal = 16'b0000001101011000;
            15'd7030: log10_cal = 16'b0000001101011000;
            15'd7031: log10_cal = 16'b0000001101011000;
            15'd7032: log10_cal = 16'b0000001101011000;
            15'd7033: log10_cal = 16'b0000001101011000;
            15'd7034: log10_cal = 16'b0000001101011000;
            15'd7035: log10_cal = 16'b0000001101011001;
            15'd7036: log10_cal = 16'b0000001101011001;
            15'd7037: log10_cal = 16'b0000001101011001;
            15'd7038: log10_cal = 16'b0000001101011001;
            15'd7039: log10_cal = 16'b0000001101011001;
            15'd7040: log10_cal = 16'b0000001101011001;
            15'd7041: log10_cal = 16'b0000001101011001;
            15'd7042: log10_cal = 16'b0000001101011001;
            15'd7043: log10_cal = 16'b0000001101011001;
            15'd7044: log10_cal = 16'b0000001101011001;
            15'd7045: log10_cal = 16'b0000001101011001;
            15'd7046: log10_cal = 16'b0000001101011001;
            15'd7047: log10_cal = 16'b0000001101011001;
            15'd7048: log10_cal = 16'b0000001101011001;
            15'd7049: log10_cal = 16'b0000001101011001;
            15'd7050: log10_cal = 16'b0000001101011001;
            15'd7051: log10_cal = 16'b0000001101011010;
            15'd7052: log10_cal = 16'b0000001101011010;
            15'd7053: log10_cal = 16'b0000001101011010;
            15'd7054: log10_cal = 16'b0000001101011010;
            15'd7055: log10_cal = 16'b0000001101011010;
            15'd7056: log10_cal = 16'b0000001101011010;
            15'd7057: log10_cal = 16'b0000001101011010;
            15'd7058: log10_cal = 16'b0000001101011010;
            15'd7059: log10_cal = 16'b0000001101011010;
            15'd7060: log10_cal = 16'b0000001101011010;
            15'd7061: log10_cal = 16'b0000001101011010;
            15'd7062: log10_cal = 16'b0000001101011010;
            15'd7063: log10_cal = 16'b0000001101011010;
            15'd7064: log10_cal = 16'b0000001101011010;
            15'd7065: log10_cal = 16'b0000001101011010;
            15'd7066: log10_cal = 16'b0000001101011011;
            15'd7067: log10_cal = 16'b0000001101011011;
            15'd7068: log10_cal = 16'b0000001101011011;
            15'd7069: log10_cal = 16'b0000001101011011;
            15'd7070: log10_cal = 16'b0000001101011011;
            15'd7071: log10_cal = 16'b0000001101011011;
            15'd7072: log10_cal = 16'b0000001101011011;
            15'd7073: log10_cal = 16'b0000001101011011;
            15'd7074: log10_cal = 16'b0000001101011011;
            15'd7075: log10_cal = 16'b0000001101011011;
            15'd7076: log10_cal = 16'b0000001101011011;
            15'd7077: log10_cal = 16'b0000001101011011;
            15'd7078: log10_cal = 16'b0000001101011011;
            15'd7079: log10_cal = 16'b0000001101011011;
            15'd7080: log10_cal = 16'b0000001101011011;
            15'd7081: log10_cal = 16'b0000001101011011;
            15'd7082: log10_cal = 16'b0000001101011100;
            15'd7083: log10_cal = 16'b0000001101011100;
            15'd7084: log10_cal = 16'b0000001101011100;
            15'd7085: log10_cal = 16'b0000001101011100;
            15'd7086: log10_cal = 16'b0000001101011100;
            15'd7087: log10_cal = 16'b0000001101011100;
            15'd7088: log10_cal = 16'b0000001101011100;
            15'd7089: log10_cal = 16'b0000001101011100;
            15'd7090: log10_cal = 16'b0000001101011100;
            15'd7091: log10_cal = 16'b0000001101011100;
            15'd7092: log10_cal = 16'b0000001101011100;
            15'd7093: log10_cal = 16'b0000001101011100;
            15'd7094: log10_cal = 16'b0000001101011100;
            15'd7095: log10_cal = 16'b0000001101011100;
            15'd7096: log10_cal = 16'b0000001101011100;
            15'd7097: log10_cal = 16'b0000001101011100;
            15'd7098: log10_cal = 16'b0000001101011101;
            15'd7099: log10_cal = 16'b0000001101011101;
            15'd7100: log10_cal = 16'b0000001101011101;
            15'd7101: log10_cal = 16'b0000001101011101;
            15'd7102: log10_cal = 16'b0000001101011101;
            15'd7103: log10_cal = 16'b0000001101011101;
            15'd7104: log10_cal = 16'b0000001101011101;
            15'd7105: log10_cal = 16'b0000001101011101;
            15'd7106: log10_cal = 16'b0000001101011101;
            15'd7107: log10_cal = 16'b0000001101011101;
            15'd7108: log10_cal = 16'b0000001101011101;
            15'd7109: log10_cal = 16'b0000001101011101;
            15'd7110: log10_cal = 16'b0000001101011101;
            15'd7111: log10_cal = 16'b0000001101011101;
            15'd7112: log10_cal = 16'b0000001101011101;
            15'd7113: log10_cal = 16'b0000001101011101;
            15'd7114: log10_cal = 16'b0000001101011110;
            15'd7115: log10_cal = 16'b0000001101011110;
            15'd7116: log10_cal = 16'b0000001101011110;
            15'd7117: log10_cal = 16'b0000001101011110;
            15'd7118: log10_cal = 16'b0000001101011110;
            15'd7119: log10_cal = 16'b0000001101011110;
            15'd7120: log10_cal = 16'b0000001101011110;
            15'd7121: log10_cal = 16'b0000001101011110;
            15'd7122: log10_cal = 16'b0000001101011110;
            15'd7123: log10_cal = 16'b0000001101011110;
            15'd7124: log10_cal = 16'b0000001101011110;
            15'd7125: log10_cal = 16'b0000001101011110;
            15'd7126: log10_cal = 16'b0000001101011110;
            15'd7127: log10_cal = 16'b0000001101011110;
            15'd7128: log10_cal = 16'b0000001101011110;
            15'd7129: log10_cal = 16'b0000001101011110;
            15'd7130: log10_cal = 16'b0000001101011111;
            15'd7131: log10_cal = 16'b0000001101011111;
            15'd7132: log10_cal = 16'b0000001101011111;
            15'd7133: log10_cal = 16'b0000001101011111;
            15'd7134: log10_cal = 16'b0000001101011111;
            15'd7135: log10_cal = 16'b0000001101011111;
            15'd7136: log10_cal = 16'b0000001101011111;
            15'd7137: log10_cal = 16'b0000001101011111;
            15'd7138: log10_cal = 16'b0000001101011111;
            15'd7139: log10_cal = 16'b0000001101011111;
            15'd7140: log10_cal = 16'b0000001101011111;
            15'd7141: log10_cal = 16'b0000001101011111;
            15'd7142: log10_cal = 16'b0000001101011111;
            15'd7143: log10_cal = 16'b0000001101011111;
            15'd7144: log10_cal = 16'b0000001101011111;
            15'd7145: log10_cal = 16'b0000001101011111;
            15'd7146: log10_cal = 16'b0000001101100000;
            15'd7147: log10_cal = 16'b0000001101100000;
            15'd7148: log10_cal = 16'b0000001101100000;
            15'd7149: log10_cal = 16'b0000001101100000;
            15'd7150: log10_cal = 16'b0000001101100000;
            15'd7151: log10_cal = 16'b0000001101100000;
            15'd7152: log10_cal = 16'b0000001101100000;
            15'd7153: log10_cal = 16'b0000001101100000;
            15'd7154: log10_cal = 16'b0000001101100000;
            15'd7155: log10_cal = 16'b0000001101100000;
            15'd7156: log10_cal = 16'b0000001101100000;
            15'd7157: log10_cal = 16'b0000001101100000;
            15'd7158: log10_cal = 16'b0000001101100000;
            15'd7159: log10_cal = 16'b0000001101100000;
            15'd7160: log10_cal = 16'b0000001101100000;
            15'd7161: log10_cal = 16'b0000001101100000;
            15'd7162: log10_cal = 16'b0000001101100001;
            15'd7163: log10_cal = 16'b0000001101100001;
            15'd7164: log10_cal = 16'b0000001101100001;
            15'd7165: log10_cal = 16'b0000001101100001;
            15'd7166: log10_cal = 16'b0000001101100001;
            15'd7167: log10_cal = 16'b0000001101100001;
            15'd7168: log10_cal = 16'b0000001101100001;
            15'd7169: log10_cal = 16'b0000001101100001;
            15'd7170: log10_cal = 16'b0000001101100001;
            15'd7171: log10_cal = 16'b0000001101100001;
            15'd7172: log10_cal = 16'b0000001101100001;
            15'd7173: log10_cal = 16'b0000001101100001;
            15'd7174: log10_cal = 16'b0000001101100001;
            15'd7175: log10_cal = 16'b0000001101100001;
            15'd7176: log10_cal = 16'b0000001101100001;
            15'd7177: log10_cal = 16'b0000001101100001;
            15'd7178: log10_cal = 16'b0000001101100010;
            15'd7179: log10_cal = 16'b0000001101100010;
            15'd7180: log10_cal = 16'b0000001101100010;
            15'd7181: log10_cal = 16'b0000001101100010;
            15'd7182: log10_cal = 16'b0000001101100010;
            15'd7183: log10_cal = 16'b0000001101100010;
            15'd7184: log10_cal = 16'b0000001101100010;
            15'd7185: log10_cal = 16'b0000001101100010;
            15'd7186: log10_cal = 16'b0000001101100010;
            15'd7187: log10_cal = 16'b0000001101100010;
            15'd7188: log10_cal = 16'b0000001101100010;
            15'd7189: log10_cal = 16'b0000001101100010;
            15'd7190: log10_cal = 16'b0000001101100010;
            15'd7191: log10_cal = 16'b0000001101100010;
            15'd7192: log10_cal = 16'b0000001101100010;
            15'd7193: log10_cal = 16'b0000001101100010;
            15'd7194: log10_cal = 16'b0000001101100010;
            15'd7195: log10_cal = 16'b0000001101100011;
            15'd7196: log10_cal = 16'b0000001101100011;
            15'd7197: log10_cal = 16'b0000001101100011;
            15'd7198: log10_cal = 16'b0000001101100011;
            15'd7199: log10_cal = 16'b0000001101100011;
            15'd7200: log10_cal = 16'b0000001101100011;
            15'd7201: log10_cal = 16'b0000001101100011;
            15'd7202: log10_cal = 16'b0000001101100011;
            15'd7203: log10_cal = 16'b0000001101100011;
            15'd7204: log10_cal = 16'b0000001101100011;
            15'd7205: log10_cal = 16'b0000001101100011;
            15'd7206: log10_cal = 16'b0000001101100011;
            15'd7207: log10_cal = 16'b0000001101100011;
            15'd7208: log10_cal = 16'b0000001101100011;
            15'd7209: log10_cal = 16'b0000001101100011;
            15'd7210: log10_cal = 16'b0000001101100011;
            15'd7211: log10_cal = 16'b0000001101100100;
            15'd7212: log10_cal = 16'b0000001101100100;
            15'd7213: log10_cal = 16'b0000001101100100;
            15'd7214: log10_cal = 16'b0000001101100100;
            15'd7215: log10_cal = 16'b0000001101100100;
            15'd7216: log10_cal = 16'b0000001101100100;
            15'd7217: log10_cal = 16'b0000001101100100;
            15'd7218: log10_cal = 16'b0000001101100100;
            15'd7219: log10_cal = 16'b0000001101100100;
            15'd7220: log10_cal = 16'b0000001101100100;
            15'd7221: log10_cal = 16'b0000001101100100;
            15'd7222: log10_cal = 16'b0000001101100100;
            15'd7223: log10_cal = 16'b0000001101100100;
            15'd7224: log10_cal = 16'b0000001101100100;
            15'd7225: log10_cal = 16'b0000001101100100;
            15'd7226: log10_cal = 16'b0000001101100100;
            15'd7227: log10_cal = 16'b0000001101100101;
            15'd7228: log10_cal = 16'b0000001101100101;
            15'd7229: log10_cal = 16'b0000001101100101;
            15'd7230: log10_cal = 16'b0000001101100101;
            15'd7231: log10_cal = 16'b0000001101100101;
            15'd7232: log10_cal = 16'b0000001101100101;
            15'd7233: log10_cal = 16'b0000001101100101;
            15'd7234: log10_cal = 16'b0000001101100101;
            15'd7235: log10_cal = 16'b0000001101100101;
            15'd7236: log10_cal = 16'b0000001101100101;
            15'd7237: log10_cal = 16'b0000001101100101;
            15'd7238: log10_cal = 16'b0000001101100101;
            15'd7239: log10_cal = 16'b0000001101100101;
            15'd7240: log10_cal = 16'b0000001101100101;
            15'd7241: log10_cal = 16'b0000001101100101;
            15'd7242: log10_cal = 16'b0000001101100101;
            15'd7243: log10_cal = 16'b0000001101100110;
            15'd7244: log10_cal = 16'b0000001101100110;
            15'd7245: log10_cal = 16'b0000001101100110;
            15'd7246: log10_cal = 16'b0000001101100110;
            15'd7247: log10_cal = 16'b0000001101100110;
            15'd7248: log10_cal = 16'b0000001101100110;
            15'd7249: log10_cal = 16'b0000001101100110;
            15'd7250: log10_cal = 16'b0000001101100110;
            15'd7251: log10_cal = 16'b0000001101100110;
            15'd7252: log10_cal = 16'b0000001101100110;
            15'd7253: log10_cal = 16'b0000001101100110;
            15'd7254: log10_cal = 16'b0000001101100110;
            15'd7255: log10_cal = 16'b0000001101100110;
            15'd7256: log10_cal = 16'b0000001101100110;
            15'd7257: log10_cal = 16'b0000001101100110;
            15'd7258: log10_cal = 16'b0000001101100110;
            15'd7259: log10_cal = 16'b0000001101100110;
            15'd7260: log10_cal = 16'b0000001101100111;
            15'd7261: log10_cal = 16'b0000001101100111;
            15'd7262: log10_cal = 16'b0000001101100111;
            15'd7263: log10_cal = 16'b0000001101100111;
            15'd7264: log10_cal = 16'b0000001101100111;
            15'd7265: log10_cal = 16'b0000001101100111;
            15'd7266: log10_cal = 16'b0000001101100111;
            15'd7267: log10_cal = 16'b0000001101100111;
            15'd7268: log10_cal = 16'b0000001101100111;
            15'd7269: log10_cal = 16'b0000001101100111;
            15'd7270: log10_cal = 16'b0000001101100111;
            15'd7271: log10_cal = 16'b0000001101100111;
            15'd7272: log10_cal = 16'b0000001101100111;
            15'd7273: log10_cal = 16'b0000001101100111;
            15'd7274: log10_cal = 16'b0000001101100111;
            15'd7275: log10_cal = 16'b0000001101100111;
            15'd7276: log10_cal = 16'b0000001101101000;
            15'd7277: log10_cal = 16'b0000001101101000;
            15'd7278: log10_cal = 16'b0000001101101000;
            15'd7279: log10_cal = 16'b0000001101101000;
            15'd7280: log10_cal = 16'b0000001101101000;
            15'd7281: log10_cal = 16'b0000001101101000;
            15'd7282: log10_cal = 16'b0000001101101000;
            15'd7283: log10_cal = 16'b0000001101101000;
            15'd7284: log10_cal = 16'b0000001101101000;
            15'd7285: log10_cal = 16'b0000001101101000;
            15'd7286: log10_cal = 16'b0000001101101000;
            15'd7287: log10_cal = 16'b0000001101101000;
            15'd7288: log10_cal = 16'b0000001101101000;
            15'd7289: log10_cal = 16'b0000001101101000;
            15'd7290: log10_cal = 16'b0000001101101000;
            15'd7291: log10_cal = 16'b0000001101101000;
            15'd7292: log10_cal = 16'b0000001101101001;
            15'd7293: log10_cal = 16'b0000001101101001;
            15'd7294: log10_cal = 16'b0000001101101001;
            15'd7295: log10_cal = 16'b0000001101101001;
            15'd7296: log10_cal = 16'b0000001101101001;
            15'd7297: log10_cal = 16'b0000001101101001;
            15'd7298: log10_cal = 16'b0000001101101001;
            15'd7299: log10_cal = 16'b0000001101101001;
            15'd7300: log10_cal = 16'b0000001101101001;
            15'd7301: log10_cal = 16'b0000001101101001;
            15'd7302: log10_cal = 16'b0000001101101001;
            15'd7303: log10_cal = 16'b0000001101101001;
            15'd7304: log10_cal = 16'b0000001101101001;
            15'd7305: log10_cal = 16'b0000001101101001;
            15'd7306: log10_cal = 16'b0000001101101001;
            15'd7307: log10_cal = 16'b0000001101101001;
            15'd7308: log10_cal = 16'b0000001101101001;
            15'd7309: log10_cal = 16'b0000001101101010;
            15'd7310: log10_cal = 16'b0000001101101010;
            15'd7311: log10_cal = 16'b0000001101101010;
            15'd7312: log10_cal = 16'b0000001101101010;
            15'd7313: log10_cal = 16'b0000001101101010;
            15'd7314: log10_cal = 16'b0000001101101010;
            15'd7315: log10_cal = 16'b0000001101101010;
            15'd7316: log10_cal = 16'b0000001101101010;
            15'd7317: log10_cal = 16'b0000001101101010;
            15'd7318: log10_cal = 16'b0000001101101010;
            15'd7319: log10_cal = 16'b0000001101101010;
            15'd7320: log10_cal = 16'b0000001101101010;
            15'd7321: log10_cal = 16'b0000001101101010;
            15'd7322: log10_cal = 16'b0000001101101010;
            15'd7323: log10_cal = 16'b0000001101101010;
            15'd7324: log10_cal = 16'b0000001101101010;
            15'd7325: log10_cal = 16'b0000001101101011;
            15'd7326: log10_cal = 16'b0000001101101011;
            15'd7327: log10_cal = 16'b0000001101101011;
            15'd7328: log10_cal = 16'b0000001101101011;
            15'd7329: log10_cal = 16'b0000001101101011;
            15'd7330: log10_cal = 16'b0000001101101011;
            15'd7331: log10_cal = 16'b0000001101101011;
            15'd7332: log10_cal = 16'b0000001101101011;
            15'd7333: log10_cal = 16'b0000001101101011;
            15'd7334: log10_cal = 16'b0000001101101011;
            15'd7335: log10_cal = 16'b0000001101101011;
            15'd7336: log10_cal = 16'b0000001101101011;
            15'd7337: log10_cal = 16'b0000001101101011;
            15'd7338: log10_cal = 16'b0000001101101011;
            15'd7339: log10_cal = 16'b0000001101101011;
            15'd7340: log10_cal = 16'b0000001101101011;
            15'd7341: log10_cal = 16'b0000001101101011;
            15'd7342: log10_cal = 16'b0000001101101100;
            15'd7343: log10_cal = 16'b0000001101101100;
            15'd7344: log10_cal = 16'b0000001101101100;
            15'd7345: log10_cal = 16'b0000001101101100;
            15'd7346: log10_cal = 16'b0000001101101100;
            15'd7347: log10_cal = 16'b0000001101101100;
            15'd7348: log10_cal = 16'b0000001101101100;
            15'd7349: log10_cal = 16'b0000001101101100;
            15'd7350: log10_cal = 16'b0000001101101100;
            15'd7351: log10_cal = 16'b0000001101101100;
            15'd7352: log10_cal = 16'b0000001101101100;
            15'd7353: log10_cal = 16'b0000001101101100;
            15'd7354: log10_cal = 16'b0000001101101100;
            15'd7355: log10_cal = 16'b0000001101101100;
            15'd7356: log10_cal = 16'b0000001101101100;
            15'd7357: log10_cal = 16'b0000001101101100;
            15'd7358: log10_cal = 16'b0000001101101101;
            15'd7359: log10_cal = 16'b0000001101101101;
            15'd7360: log10_cal = 16'b0000001101101101;
            15'd7361: log10_cal = 16'b0000001101101101;
            15'd7362: log10_cal = 16'b0000001101101101;
            15'd7363: log10_cal = 16'b0000001101101101;
            15'd7364: log10_cal = 16'b0000001101101101;
            15'd7365: log10_cal = 16'b0000001101101101;
            15'd7366: log10_cal = 16'b0000001101101101;
            15'd7367: log10_cal = 16'b0000001101101101;
            15'd7368: log10_cal = 16'b0000001101101101;
            15'd7369: log10_cal = 16'b0000001101101101;
            15'd7370: log10_cal = 16'b0000001101101101;
            15'd7371: log10_cal = 16'b0000001101101101;
            15'd7372: log10_cal = 16'b0000001101101101;
            15'd7373: log10_cal = 16'b0000001101101101;
            15'd7374: log10_cal = 16'b0000001101101101;
            15'd7375: log10_cal = 16'b0000001101101110;
            15'd7376: log10_cal = 16'b0000001101101110;
            15'd7377: log10_cal = 16'b0000001101101110;
            15'd7378: log10_cal = 16'b0000001101101110;
            15'd7379: log10_cal = 16'b0000001101101110;
            15'd7380: log10_cal = 16'b0000001101101110;
            15'd7381: log10_cal = 16'b0000001101101110;
            15'd7382: log10_cal = 16'b0000001101101110;
            15'd7383: log10_cal = 16'b0000001101101110;
            15'd7384: log10_cal = 16'b0000001101101110;
            15'd7385: log10_cal = 16'b0000001101101110;
            15'd7386: log10_cal = 16'b0000001101101110;
            15'd7387: log10_cal = 16'b0000001101101110;
            15'd7388: log10_cal = 16'b0000001101101110;
            15'd7389: log10_cal = 16'b0000001101101110;
            15'd7390: log10_cal = 16'b0000001101101110;
            15'd7391: log10_cal = 16'b0000001101101111;
            15'd7392: log10_cal = 16'b0000001101101111;
            15'd7393: log10_cal = 16'b0000001101101111;
            15'd7394: log10_cal = 16'b0000001101101111;
            15'd7395: log10_cal = 16'b0000001101101111;
            15'd7396: log10_cal = 16'b0000001101101111;
            15'd7397: log10_cal = 16'b0000001101101111;
            15'd7398: log10_cal = 16'b0000001101101111;
            15'd7399: log10_cal = 16'b0000001101101111;
            15'd7400: log10_cal = 16'b0000001101101111;
            15'd7401: log10_cal = 16'b0000001101101111;
            15'd7402: log10_cal = 16'b0000001101101111;
            15'd7403: log10_cal = 16'b0000001101101111;
            15'd7404: log10_cal = 16'b0000001101101111;
            15'd7405: log10_cal = 16'b0000001101101111;
            15'd7406: log10_cal = 16'b0000001101101111;
            15'd7407: log10_cal = 16'b0000001101101111;
            15'd7408: log10_cal = 16'b0000001101110000;
            15'd7409: log10_cal = 16'b0000001101110000;
            15'd7410: log10_cal = 16'b0000001101110000;
            15'd7411: log10_cal = 16'b0000001101110000;
            15'd7412: log10_cal = 16'b0000001101110000;
            15'd7413: log10_cal = 16'b0000001101110000;
            15'd7414: log10_cal = 16'b0000001101110000;
            15'd7415: log10_cal = 16'b0000001101110000;
            15'd7416: log10_cal = 16'b0000001101110000;
            15'd7417: log10_cal = 16'b0000001101110000;
            15'd7418: log10_cal = 16'b0000001101110000;
            15'd7419: log10_cal = 16'b0000001101110000;
            15'd7420: log10_cal = 16'b0000001101110000;
            15'd7421: log10_cal = 16'b0000001101110000;
            15'd7422: log10_cal = 16'b0000001101110000;
            15'd7423: log10_cal = 16'b0000001101110000;
            15'd7424: log10_cal = 16'b0000001101110000;
            15'd7425: log10_cal = 16'b0000001101110001;
            15'd7426: log10_cal = 16'b0000001101110001;
            15'd7427: log10_cal = 16'b0000001101110001;
            15'd7428: log10_cal = 16'b0000001101110001;
            15'd7429: log10_cal = 16'b0000001101110001;
            15'd7430: log10_cal = 16'b0000001101110001;
            15'd7431: log10_cal = 16'b0000001101110001;
            15'd7432: log10_cal = 16'b0000001101110001;
            15'd7433: log10_cal = 16'b0000001101110001;
            15'd7434: log10_cal = 16'b0000001101110001;
            15'd7435: log10_cal = 16'b0000001101110001;
            15'd7436: log10_cal = 16'b0000001101110001;
            15'd7437: log10_cal = 16'b0000001101110001;
            15'd7438: log10_cal = 16'b0000001101110001;
            15'd7439: log10_cal = 16'b0000001101110001;
            15'd7440: log10_cal = 16'b0000001101110001;
            15'd7441: log10_cal = 16'b0000001101110010;
            15'd7442: log10_cal = 16'b0000001101110010;
            15'd7443: log10_cal = 16'b0000001101110010;
            15'd7444: log10_cal = 16'b0000001101110010;
            15'd7445: log10_cal = 16'b0000001101110010;
            15'd7446: log10_cal = 16'b0000001101110010;
            15'd7447: log10_cal = 16'b0000001101110010;
            15'd7448: log10_cal = 16'b0000001101110010;
            15'd7449: log10_cal = 16'b0000001101110010;
            15'd7450: log10_cal = 16'b0000001101110010;
            15'd7451: log10_cal = 16'b0000001101110010;
            15'd7452: log10_cal = 16'b0000001101110010;
            15'd7453: log10_cal = 16'b0000001101110010;
            15'd7454: log10_cal = 16'b0000001101110010;
            15'd7455: log10_cal = 16'b0000001101110010;
            15'd7456: log10_cal = 16'b0000001101110010;
            15'd7457: log10_cal = 16'b0000001101110010;
            15'd7458: log10_cal = 16'b0000001101110011;
            15'd7459: log10_cal = 16'b0000001101110011;
            15'd7460: log10_cal = 16'b0000001101110011;
            15'd7461: log10_cal = 16'b0000001101110011;
            15'd7462: log10_cal = 16'b0000001101110011;
            15'd7463: log10_cal = 16'b0000001101110011;
            15'd7464: log10_cal = 16'b0000001101110011;
            15'd7465: log10_cal = 16'b0000001101110011;
            15'd7466: log10_cal = 16'b0000001101110011;
            15'd7467: log10_cal = 16'b0000001101110011;
            15'd7468: log10_cal = 16'b0000001101110011;
            15'd7469: log10_cal = 16'b0000001101110011;
            15'd7470: log10_cal = 16'b0000001101110011;
            15'd7471: log10_cal = 16'b0000001101110011;
            15'd7472: log10_cal = 16'b0000001101110011;
            15'd7473: log10_cal = 16'b0000001101110011;
            15'd7474: log10_cal = 16'b0000001101110011;
            15'd7475: log10_cal = 16'b0000001101110100;
            15'd7476: log10_cal = 16'b0000001101110100;
            15'd7477: log10_cal = 16'b0000001101110100;
            15'd7478: log10_cal = 16'b0000001101110100;
            15'd7479: log10_cal = 16'b0000001101110100;
            15'd7480: log10_cal = 16'b0000001101110100;
            15'd7481: log10_cal = 16'b0000001101110100;
            15'd7482: log10_cal = 16'b0000001101110100;
            15'd7483: log10_cal = 16'b0000001101110100;
            15'd7484: log10_cal = 16'b0000001101110100;
            15'd7485: log10_cal = 16'b0000001101110100;
            15'd7486: log10_cal = 16'b0000001101110100;
            15'd7487: log10_cal = 16'b0000001101110100;
            15'd7488: log10_cal = 16'b0000001101110100;
            15'd7489: log10_cal = 16'b0000001101110100;
            15'd7490: log10_cal = 16'b0000001101110100;
            15'd7491: log10_cal = 16'b0000001101110100;
            15'd7492: log10_cal = 16'b0000001101110101;
            15'd7493: log10_cal = 16'b0000001101110101;
            15'd7494: log10_cal = 16'b0000001101110101;
            15'd7495: log10_cal = 16'b0000001101110101;
            15'd7496: log10_cal = 16'b0000001101110101;
            15'd7497: log10_cal = 16'b0000001101110101;
            15'd7498: log10_cal = 16'b0000001101110101;
            15'd7499: log10_cal = 16'b0000001101110101;
            15'd7500: log10_cal = 16'b0000001101110101;
            15'd7501: log10_cal = 16'b0000001101110101;
            15'd7502: log10_cal = 16'b0000001101110101;
            15'd7503: log10_cal = 16'b0000001101110101;
            15'd7504: log10_cal = 16'b0000001101110101;
            15'd7505: log10_cal = 16'b0000001101110101;
            15'd7506: log10_cal = 16'b0000001101110101;
            15'd7507: log10_cal = 16'b0000001101110101;
            15'd7508: log10_cal = 16'b0000001101110101;
            15'd7509: log10_cal = 16'b0000001101110110;
            15'd7510: log10_cal = 16'b0000001101110110;
            15'd7511: log10_cal = 16'b0000001101110110;
            15'd7512: log10_cal = 16'b0000001101110110;
            15'd7513: log10_cal = 16'b0000001101110110;
            15'd7514: log10_cal = 16'b0000001101110110;
            15'd7515: log10_cal = 16'b0000001101110110;
            15'd7516: log10_cal = 16'b0000001101110110;
            15'd7517: log10_cal = 16'b0000001101110110;
            15'd7518: log10_cal = 16'b0000001101110110;
            15'd7519: log10_cal = 16'b0000001101110110;
            15'd7520: log10_cal = 16'b0000001101110110;
            15'd7521: log10_cal = 16'b0000001101110110;
            15'd7522: log10_cal = 16'b0000001101110110;
            15'd7523: log10_cal = 16'b0000001101110110;
            15'd7524: log10_cal = 16'b0000001101110110;
            15'd7525: log10_cal = 16'b0000001101110110;
            15'd7526: log10_cal = 16'b0000001101110111;
            15'd7527: log10_cal = 16'b0000001101110111;
            15'd7528: log10_cal = 16'b0000001101110111;
            15'd7529: log10_cal = 16'b0000001101110111;
            15'd7530: log10_cal = 16'b0000001101110111;
            15'd7531: log10_cal = 16'b0000001101110111;
            15'd7532: log10_cal = 16'b0000001101110111;
            15'd7533: log10_cal = 16'b0000001101110111;
            15'd7534: log10_cal = 16'b0000001101110111;
            15'd7535: log10_cal = 16'b0000001101110111;
            15'd7536: log10_cal = 16'b0000001101110111;
            15'd7537: log10_cal = 16'b0000001101110111;
            15'd7538: log10_cal = 16'b0000001101110111;
            15'd7539: log10_cal = 16'b0000001101110111;
            15'd7540: log10_cal = 16'b0000001101110111;
            15'd7541: log10_cal = 16'b0000001101110111;
            15'd7542: log10_cal = 16'b0000001101110111;
            15'd7543: log10_cal = 16'b0000001101111000;
            15'd7544: log10_cal = 16'b0000001101111000;
            15'd7545: log10_cal = 16'b0000001101111000;
            15'd7546: log10_cal = 16'b0000001101111000;
            15'd7547: log10_cal = 16'b0000001101111000;
            15'd7548: log10_cal = 16'b0000001101111000;
            15'd7549: log10_cal = 16'b0000001101111000;
            15'd7550: log10_cal = 16'b0000001101111000;
            15'd7551: log10_cal = 16'b0000001101111000;
            15'd7552: log10_cal = 16'b0000001101111000;
            15'd7553: log10_cal = 16'b0000001101111000;
            15'd7554: log10_cal = 16'b0000001101111000;
            15'd7555: log10_cal = 16'b0000001101111000;
            15'd7556: log10_cal = 16'b0000001101111000;
            15'd7557: log10_cal = 16'b0000001101111000;
            15'd7558: log10_cal = 16'b0000001101111000;
            15'd7559: log10_cal = 16'b0000001101111001;
            15'd7560: log10_cal = 16'b0000001101111001;
            15'd7561: log10_cal = 16'b0000001101111001;
            15'd7562: log10_cal = 16'b0000001101111001;
            15'd7563: log10_cal = 16'b0000001101111001;
            15'd7564: log10_cal = 16'b0000001101111001;
            15'd7565: log10_cal = 16'b0000001101111001;
            15'd7566: log10_cal = 16'b0000001101111001;
            15'd7567: log10_cal = 16'b0000001101111001;
            15'd7568: log10_cal = 16'b0000001101111001;
            15'd7569: log10_cal = 16'b0000001101111001;
            15'd7570: log10_cal = 16'b0000001101111001;
            15'd7571: log10_cal = 16'b0000001101111001;
            15'd7572: log10_cal = 16'b0000001101111001;
            15'd7573: log10_cal = 16'b0000001101111001;
            15'd7574: log10_cal = 16'b0000001101111001;
            15'd7575: log10_cal = 16'b0000001101111001;
            15'd7576: log10_cal = 16'b0000001101111001;
            15'd7577: log10_cal = 16'b0000001101111010;
            15'd7578: log10_cal = 16'b0000001101111010;
            15'd7579: log10_cal = 16'b0000001101111010;
            15'd7580: log10_cal = 16'b0000001101111010;
            15'd7581: log10_cal = 16'b0000001101111010;
            15'd7582: log10_cal = 16'b0000001101111010;
            15'd7583: log10_cal = 16'b0000001101111010;
            15'd7584: log10_cal = 16'b0000001101111010;
            15'd7585: log10_cal = 16'b0000001101111010;
            15'd7586: log10_cal = 16'b0000001101111010;
            15'd7587: log10_cal = 16'b0000001101111010;
            15'd7588: log10_cal = 16'b0000001101111010;
            15'd7589: log10_cal = 16'b0000001101111010;
            15'd7590: log10_cal = 16'b0000001101111010;
            15'd7591: log10_cal = 16'b0000001101111010;
            15'd7592: log10_cal = 16'b0000001101111010;
            15'd7593: log10_cal = 16'b0000001101111010;
            15'd7594: log10_cal = 16'b0000001101111011;
            15'd7595: log10_cal = 16'b0000001101111011;
            15'd7596: log10_cal = 16'b0000001101111011;
            15'd7597: log10_cal = 16'b0000001101111011;
            15'd7598: log10_cal = 16'b0000001101111011;
            15'd7599: log10_cal = 16'b0000001101111011;
            15'd7600: log10_cal = 16'b0000001101111011;
            15'd7601: log10_cal = 16'b0000001101111011;
            15'd7602: log10_cal = 16'b0000001101111011;
            15'd7603: log10_cal = 16'b0000001101111011;
            15'd7604: log10_cal = 16'b0000001101111011;
            15'd7605: log10_cal = 16'b0000001101111011;
            15'd7606: log10_cal = 16'b0000001101111011;
            15'd7607: log10_cal = 16'b0000001101111011;
            15'd7608: log10_cal = 16'b0000001101111011;
            15'd7609: log10_cal = 16'b0000001101111011;
            15'd7610: log10_cal = 16'b0000001101111011;
            15'd7611: log10_cal = 16'b0000001101111100;
            15'd7612: log10_cal = 16'b0000001101111100;
            15'd7613: log10_cal = 16'b0000001101111100;
            15'd7614: log10_cal = 16'b0000001101111100;
            15'd7615: log10_cal = 16'b0000001101111100;
            15'd7616: log10_cal = 16'b0000001101111100;
            15'd7617: log10_cal = 16'b0000001101111100;
            15'd7618: log10_cal = 16'b0000001101111100;
            15'd7619: log10_cal = 16'b0000001101111100;
            15'd7620: log10_cal = 16'b0000001101111100;
            15'd7621: log10_cal = 16'b0000001101111100;
            15'd7622: log10_cal = 16'b0000001101111100;
            15'd7623: log10_cal = 16'b0000001101111100;
            15'd7624: log10_cal = 16'b0000001101111100;
            15'd7625: log10_cal = 16'b0000001101111100;
            15'd7626: log10_cal = 16'b0000001101111100;
            15'd7627: log10_cal = 16'b0000001101111100;
            15'd7628: log10_cal = 16'b0000001101111101;
            15'd7629: log10_cal = 16'b0000001101111101;
            15'd7630: log10_cal = 16'b0000001101111101;
            15'd7631: log10_cal = 16'b0000001101111101;
            15'd7632: log10_cal = 16'b0000001101111101;
            15'd7633: log10_cal = 16'b0000001101111101;
            15'd7634: log10_cal = 16'b0000001101111101;
            15'd7635: log10_cal = 16'b0000001101111101;
            15'd7636: log10_cal = 16'b0000001101111101;
            15'd7637: log10_cal = 16'b0000001101111101;
            15'd7638: log10_cal = 16'b0000001101111101;
            15'd7639: log10_cal = 16'b0000001101111101;
            15'd7640: log10_cal = 16'b0000001101111101;
            15'd7641: log10_cal = 16'b0000001101111101;
            15'd7642: log10_cal = 16'b0000001101111101;
            15'd7643: log10_cal = 16'b0000001101111101;
            15'd7644: log10_cal = 16'b0000001101111101;
            15'd7645: log10_cal = 16'b0000001101111110;
            15'd7646: log10_cal = 16'b0000001101111110;
            15'd7647: log10_cal = 16'b0000001101111110;
            15'd7648: log10_cal = 16'b0000001101111110;
            15'd7649: log10_cal = 16'b0000001101111110;
            15'd7650: log10_cal = 16'b0000001101111110;
            15'd7651: log10_cal = 16'b0000001101111110;
            15'd7652: log10_cal = 16'b0000001101111110;
            15'd7653: log10_cal = 16'b0000001101111110;
            15'd7654: log10_cal = 16'b0000001101111110;
            15'd7655: log10_cal = 16'b0000001101111110;
            15'd7656: log10_cal = 16'b0000001101111110;
            15'd7657: log10_cal = 16'b0000001101111110;
            15'd7658: log10_cal = 16'b0000001101111110;
            15'd7659: log10_cal = 16'b0000001101111110;
            15'd7660: log10_cal = 16'b0000001101111110;
            15'd7661: log10_cal = 16'b0000001101111110;
            15'd7662: log10_cal = 16'b0000001101111111;
            15'd7663: log10_cal = 16'b0000001101111111;
            15'd7664: log10_cal = 16'b0000001101111111;
            15'd7665: log10_cal = 16'b0000001101111111;
            15'd7666: log10_cal = 16'b0000001101111111;
            15'd7667: log10_cal = 16'b0000001101111111;
            15'd7668: log10_cal = 16'b0000001101111111;
            15'd7669: log10_cal = 16'b0000001101111111;
            15'd7670: log10_cal = 16'b0000001101111111;
            15'd7671: log10_cal = 16'b0000001101111111;
            15'd7672: log10_cal = 16'b0000001101111111;
            15'd7673: log10_cal = 16'b0000001101111111;
            15'd7674: log10_cal = 16'b0000001101111111;
            15'd7675: log10_cal = 16'b0000001101111111;
            15'd7676: log10_cal = 16'b0000001101111111;
            15'd7677: log10_cal = 16'b0000001101111111;
            15'd7678: log10_cal = 16'b0000001101111111;
            15'd7679: log10_cal = 16'b0000001110000000;
            15'd7680: log10_cal = 16'b0000001110000000;
            15'd7681: log10_cal = 16'b0000001110000000;
            15'd7682: log10_cal = 16'b0000001110000000;
            15'd7683: log10_cal = 16'b0000001110000000;
            15'd7684: log10_cal = 16'b0000001110000000;
            15'd7685: log10_cal = 16'b0000001110000000;
            15'd7686: log10_cal = 16'b0000001110000000;
            15'd7687: log10_cal = 16'b0000001110000000;
            15'd7688: log10_cal = 16'b0000001110000000;
            15'd7689: log10_cal = 16'b0000001110000000;
            15'd7690: log10_cal = 16'b0000001110000000;
            15'd7691: log10_cal = 16'b0000001110000000;
            15'd7692: log10_cal = 16'b0000001110000000;
            15'd7693: log10_cal = 16'b0000001110000000;
            15'd7694: log10_cal = 16'b0000001110000000;
            15'd7695: log10_cal = 16'b0000001110000000;
            15'd7696: log10_cal = 16'b0000001110000000;
            15'd7697: log10_cal = 16'b0000001110000001;
            15'd7698: log10_cal = 16'b0000001110000001;
            15'd7699: log10_cal = 16'b0000001110000001;
            15'd7700: log10_cal = 16'b0000001110000001;
            15'd7701: log10_cal = 16'b0000001110000001;
            15'd7702: log10_cal = 16'b0000001110000001;
            15'd7703: log10_cal = 16'b0000001110000001;
            15'd7704: log10_cal = 16'b0000001110000001;
            15'd7705: log10_cal = 16'b0000001110000001;
            15'd7706: log10_cal = 16'b0000001110000001;
            15'd7707: log10_cal = 16'b0000001110000001;
            15'd7708: log10_cal = 16'b0000001110000001;
            15'd7709: log10_cal = 16'b0000001110000001;
            15'd7710: log10_cal = 16'b0000001110000001;
            15'd7711: log10_cal = 16'b0000001110000001;
            15'd7712: log10_cal = 16'b0000001110000001;
            15'd7713: log10_cal = 16'b0000001110000001;
            15'd7714: log10_cal = 16'b0000001110000010;
            15'd7715: log10_cal = 16'b0000001110000010;
            15'd7716: log10_cal = 16'b0000001110000010;
            15'd7717: log10_cal = 16'b0000001110000010;
            15'd7718: log10_cal = 16'b0000001110000010;
            15'd7719: log10_cal = 16'b0000001110000010;
            15'd7720: log10_cal = 16'b0000001110000010;
            15'd7721: log10_cal = 16'b0000001110000010;
            15'd7722: log10_cal = 16'b0000001110000010;
            15'd7723: log10_cal = 16'b0000001110000010;
            15'd7724: log10_cal = 16'b0000001110000010;
            15'd7725: log10_cal = 16'b0000001110000010;
            15'd7726: log10_cal = 16'b0000001110000010;
            15'd7727: log10_cal = 16'b0000001110000010;
            15'd7728: log10_cal = 16'b0000001110000010;
            15'd7729: log10_cal = 16'b0000001110000010;
            15'd7730: log10_cal = 16'b0000001110000010;
            15'd7731: log10_cal = 16'b0000001110000011;
            15'd7732: log10_cal = 16'b0000001110000011;
            15'd7733: log10_cal = 16'b0000001110000011;
            15'd7734: log10_cal = 16'b0000001110000011;
            15'd7735: log10_cal = 16'b0000001110000011;
            15'd7736: log10_cal = 16'b0000001110000011;
            15'd7737: log10_cal = 16'b0000001110000011;
            15'd7738: log10_cal = 16'b0000001110000011;
            15'd7739: log10_cal = 16'b0000001110000011;
            15'd7740: log10_cal = 16'b0000001110000011;
            15'd7741: log10_cal = 16'b0000001110000011;
            15'd7742: log10_cal = 16'b0000001110000011;
            15'd7743: log10_cal = 16'b0000001110000011;
            15'd7744: log10_cal = 16'b0000001110000011;
            15'd7745: log10_cal = 16'b0000001110000011;
            15'd7746: log10_cal = 16'b0000001110000011;
            15'd7747: log10_cal = 16'b0000001110000011;
            15'd7748: log10_cal = 16'b0000001110000011;
            15'd7749: log10_cal = 16'b0000001110000100;
            15'd7750: log10_cal = 16'b0000001110000100;
            15'd7751: log10_cal = 16'b0000001110000100;
            15'd7752: log10_cal = 16'b0000001110000100;
            15'd7753: log10_cal = 16'b0000001110000100;
            15'd7754: log10_cal = 16'b0000001110000100;
            15'd7755: log10_cal = 16'b0000001110000100;
            15'd7756: log10_cal = 16'b0000001110000100;
            15'd7757: log10_cal = 16'b0000001110000100;
            15'd7758: log10_cal = 16'b0000001110000100;
            15'd7759: log10_cal = 16'b0000001110000100;
            15'd7760: log10_cal = 16'b0000001110000100;
            15'd7761: log10_cal = 16'b0000001110000100;
            15'd7762: log10_cal = 16'b0000001110000100;
            15'd7763: log10_cal = 16'b0000001110000100;
            15'd7764: log10_cal = 16'b0000001110000100;
            15'd7765: log10_cal = 16'b0000001110000100;
            15'd7766: log10_cal = 16'b0000001110000101;
            15'd7767: log10_cal = 16'b0000001110000101;
            15'd7768: log10_cal = 16'b0000001110000101;
            15'd7769: log10_cal = 16'b0000001110000101;
            15'd7770: log10_cal = 16'b0000001110000101;
            15'd7771: log10_cal = 16'b0000001110000101;
            15'd7772: log10_cal = 16'b0000001110000101;
            15'd7773: log10_cal = 16'b0000001110000101;
            15'd7774: log10_cal = 16'b0000001110000101;
            15'd7775: log10_cal = 16'b0000001110000101;
            15'd7776: log10_cal = 16'b0000001110000101;
            15'd7777: log10_cal = 16'b0000001110000101;
            15'd7778: log10_cal = 16'b0000001110000101;
            15'd7779: log10_cal = 16'b0000001110000101;
            15'd7780: log10_cal = 16'b0000001110000101;
            15'd7781: log10_cal = 16'b0000001110000101;
            15'd7782: log10_cal = 16'b0000001110000101;
            15'd7783: log10_cal = 16'b0000001110000101;
            15'd7784: log10_cal = 16'b0000001110000110;
            15'd7785: log10_cal = 16'b0000001110000110;
            15'd7786: log10_cal = 16'b0000001110000110;
            15'd7787: log10_cal = 16'b0000001110000110;
            15'd7788: log10_cal = 16'b0000001110000110;
            15'd7789: log10_cal = 16'b0000001110000110;
            15'd7790: log10_cal = 16'b0000001110000110;
            15'd7791: log10_cal = 16'b0000001110000110;
            15'd7792: log10_cal = 16'b0000001110000110;
            15'd7793: log10_cal = 16'b0000001110000110;
            15'd7794: log10_cal = 16'b0000001110000110;
            15'd7795: log10_cal = 16'b0000001110000110;
            15'd7796: log10_cal = 16'b0000001110000110;
            15'd7797: log10_cal = 16'b0000001110000110;
            15'd7798: log10_cal = 16'b0000001110000110;
            15'd7799: log10_cal = 16'b0000001110000110;
            15'd7800: log10_cal = 16'b0000001110000110;
            15'd7801: log10_cal = 16'b0000001110000111;
            15'd7802: log10_cal = 16'b0000001110000111;
            15'd7803: log10_cal = 16'b0000001110000111;
            15'd7804: log10_cal = 16'b0000001110000111;
            15'd7805: log10_cal = 16'b0000001110000111;
            15'd7806: log10_cal = 16'b0000001110000111;
            15'd7807: log10_cal = 16'b0000001110000111;
            15'd7808: log10_cal = 16'b0000001110000111;
            15'd7809: log10_cal = 16'b0000001110000111;
            15'd7810: log10_cal = 16'b0000001110000111;
            15'd7811: log10_cal = 16'b0000001110000111;
            15'd7812: log10_cal = 16'b0000001110000111;
            15'd7813: log10_cal = 16'b0000001110000111;
            15'd7814: log10_cal = 16'b0000001110000111;
            15'd7815: log10_cal = 16'b0000001110000111;
            15'd7816: log10_cal = 16'b0000001110000111;
            15'd7817: log10_cal = 16'b0000001110000111;
            15'd7818: log10_cal = 16'b0000001110000111;
            15'd7819: log10_cal = 16'b0000001110001000;
            15'd7820: log10_cal = 16'b0000001110001000;
            15'd7821: log10_cal = 16'b0000001110001000;
            15'd7822: log10_cal = 16'b0000001110001000;
            15'd7823: log10_cal = 16'b0000001110001000;
            15'd7824: log10_cal = 16'b0000001110001000;
            15'd7825: log10_cal = 16'b0000001110001000;
            15'd7826: log10_cal = 16'b0000001110001000;
            15'd7827: log10_cal = 16'b0000001110001000;
            15'd7828: log10_cal = 16'b0000001110001000;
            15'd7829: log10_cal = 16'b0000001110001000;
            15'd7830: log10_cal = 16'b0000001110001000;
            15'd7831: log10_cal = 16'b0000001110001000;
            15'd7832: log10_cal = 16'b0000001110001000;
            15'd7833: log10_cal = 16'b0000001110001000;
            15'd7834: log10_cal = 16'b0000001110001000;
            15'd7835: log10_cal = 16'b0000001110001000;
            15'd7836: log10_cal = 16'b0000001110001001;
            15'd7837: log10_cal = 16'b0000001110001001;
            15'd7838: log10_cal = 16'b0000001110001001;
            15'd7839: log10_cal = 16'b0000001110001001;
            15'd7840: log10_cal = 16'b0000001110001001;
            15'd7841: log10_cal = 16'b0000001110001001;
            15'd7842: log10_cal = 16'b0000001110001001;
            15'd7843: log10_cal = 16'b0000001110001001;
            15'd7844: log10_cal = 16'b0000001110001001;
            15'd7845: log10_cal = 16'b0000001110001001;
            15'd7846: log10_cal = 16'b0000001110001001;
            15'd7847: log10_cal = 16'b0000001110001001;
            15'd7848: log10_cal = 16'b0000001110001001;
            15'd7849: log10_cal = 16'b0000001110001001;
            15'd7850: log10_cal = 16'b0000001110001001;
            15'd7851: log10_cal = 16'b0000001110001001;
            15'd7852: log10_cal = 16'b0000001110001001;
            15'd7853: log10_cal = 16'b0000001110001001;
            15'd7854: log10_cal = 16'b0000001110001010;
            15'd7855: log10_cal = 16'b0000001110001010;
            15'd7856: log10_cal = 16'b0000001110001010;
            15'd7857: log10_cal = 16'b0000001110001010;
            15'd7858: log10_cal = 16'b0000001110001010;
            15'd7859: log10_cal = 16'b0000001110001010;
            15'd7860: log10_cal = 16'b0000001110001010;
            15'd7861: log10_cal = 16'b0000001110001010;
            15'd7862: log10_cal = 16'b0000001110001010;
            15'd7863: log10_cal = 16'b0000001110001010;
            15'd7864: log10_cal = 16'b0000001110001010;
            15'd7865: log10_cal = 16'b0000001110001010;
            15'd7866: log10_cal = 16'b0000001110001010;
            15'd7867: log10_cal = 16'b0000001110001010;
            15'd7868: log10_cal = 16'b0000001110001010;
            15'd7869: log10_cal = 16'b0000001110001010;
            15'd7870: log10_cal = 16'b0000001110001010;
            15'd7871: log10_cal = 16'b0000001110001010;
            15'd7872: log10_cal = 16'b0000001110001011;
            15'd7873: log10_cal = 16'b0000001110001011;
            15'd7874: log10_cal = 16'b0000001110001011;
            15'd7875: log10_cal = 16'b0000001110001011;
            15'd7876: log10_cal = 16'b0000001110001011;
            15'd7877: log10_cal = 16'b0000001110001011;
            15'd7878: log10_cal = 16'b0000001110001011;
            15'd7879: log10_cal = 16'b0000001110001011;
            15'd7880: log10_cal = 16'b0000001110001011;
            15'd7881: log10_cal = 16'b0000001110001011;
            15'd7882: log10_cal = 16'b0000001110001011;
            15'd7883: log10_cal = 16'b0000001110001011;
            15'd7884: log10_cal = 16'b0000001110001011;
            15'd7885: log10_cal = 16'b0000001110001011;
            15'd7886: log10_cal = 16'b0000001110001011;
            15'd7887: log10_cal = 16'b0000001110001011;
            15'd7888: log10_cal = 16'b0000001110001011;
            15'd7889: log10_cal = 16'b0000001110001100;
            15'd7890: log10_cal = 16'b0000001110001100;
            15'd7891: log10_cal = 16'b0000001110001100;
            15'd7892: log10_cal = 16'b0000001110001100;
            15'd7893: log10_cal = 16'b0000001110001100;
            15'd7894: log10_cal = 16'b0000001110001100;
            15'd7895: log10_cal = 16'b0000001110001100;
            15'd7896: log10_cal = 16'b0000001110001100;
            15'd7897: log10_cal = 16'b0000001110001100;
            15'd7898: log10_cal = 16'b0000001110001100;
            15'd7899: log10_cal = 16'b0000001110001100;
            15'd7900: log10_cal = 16'b0000001110001100;
            15'd7901: log10_cal = 16'b0000001110001100;
            15'd7902: log10_cal = 16'b0000001110001100;
            15'd7903: log10_cal = 16'b0000001110001100;
            15'd7904: log10_cal = 16'b0000001110001100;
            15'd7905: log10_cal = 16'b0000001110001100;
            15'd7906: log10_cal = 16'b0000001110001100;
            15'd7907: log10_cal = 16'b0000001110001101;
            15'd7908: log10_cal = 16'b0000001110001101;
            15'd7909: log10_cal = 16'b0000001110001101;
            15'd7910: log10_cal = 16'b0000001110001101;
            15'd7911: log10_cal = 16'b0000001110001101;
            15'd7912: log10_cal = 16'b0000001110001101;
            15'd7913: log10_cal = 16'b0000001110001101;
            15'd7914: log10_cal = 16'b0000001110001101;
            15'd7915: log10_cal = 16'b0000001110001101;
            15'd7916: log10_cal = 16'b0000001110001101;
            15'd7917: log10_cal = 16'b0000001110001101;
            15'd7918: log10_cal = 16'b0000001110001101;
            15'd7919: log10_cal = 16'b0000001110001101;
            15'd7920: log10_cal = 16'b0000001110001101;
            15'd7921: log10_cal = 16'b0000001110001101;
            15'd7922: log10_cal = 16'b0000001110001101;
            15'd7923: log10_cal = 16'b0000001110001101;
            15'd7924: log10_cal = 16'b0000001110001101;
            15'd7925: log10_cal = 16'b0000001110001110;
            15'd7926: log10_cal = 16'b0000001110001110;
            15'd7927: log10_cal = 16'b0000001110001110;
            15'd7928: log10_cal = 16'b0000001110001110;
            15'd7929: log10_cal = 16'b0000001110001110;
            15'd7930: log10_cal = 16'b0000001110001110;
            15'd7931: log10_cal = 16'b0000001110001110;
            15'd7932: log10_cal = 16'b0000001110001110;
            15'd7933: log10_cal = 16'b0000001110001110;
            15'd7934: log10_cal = 16'b0000001110001110;
            15'd7935: log10_cal = 16'b0000001110001110;
            15'd7936: log10_cal = 16'b0000001110001110;
            15'd7937: log10_cal = 16'b0000001110001110;
            15'd7938: log10_cal = 16'b0000001110001110;
            15'd7939: log10_cal = 16'b0000001110001110;
            15'd7940: log10_cal = 16'b0000001110001110;
            15'd7941: log10_cal = 16'b0000001110001110;
            15'd7942: log10_cal = 16'b0000001110001110;
            15'd7943: log10_cal = 16'b0000001110001111;
            15'd7944: log10_cal = 16'b0000001110001111;
            15'd7945: log10_cal = 16'b0000001110001111;
            15'd7946: log10_cal = 16'b0000001110001111;
            15'd7947: log10_cal = 16'b0000001110001111;
            15'd7948: log10_cal = 16'b0000001110001111;
            15'd7949: log10_cal = 16'b0000001110001111;
            15'd7950: log10_cal = 16'b0000001110001111;
            15'd7951: log10_cal = 16'b0000001110001111;
            15'd7952: log10_cal = 16'b0000001110001111;
            15'd7953: log10_cal = 16'b0000001110001111;
            15'd7954: log10_cal = 16'b0000001110001111;
            15'd7955: log10_cal = 16'b0000001110001111;
            15'd7956: log10_cal = 16'b0000001110001111;
            15'd7957: log10_cal = 16'b0000001110001111;
            15'd7958: log10_cal = 16'b0000001110001111;
            15'd7959: log10_cal = 16'b0000001110001111;
            15'd7960: log10_cal = 16'b0000001110001111;
            15'd7961: log10_cal = 16'b0000001110010000;
            15'd7962: log10_cal = 16'b0000001110010000;
            15'd7963: log10_cal = 16'b0000001110010000;
            15'd7964: log10_cal = 16'b0000001110010000;
            15'd7965: log10_cal = 16'b0000001110010000;
            15'd7966: log10_cal = 16'b0000001110010000;
            15'd7967: log10_cal = 16'b0000001110010000;
            15'd7968: log10_cal = 16'b0000001110010000;
            15'd7969: log10_cal = 16'b0000001110010000;
            15'd7970: log10_cal = 16'b0000001110010000;
            15'd7971: log10_cal = 16'b0000001110010000;
            15'd7972: log10_cal = 16'b0000001110010000;
            15'd7973: log10_cal = 16'b0000001110010000;
            15'd7974: log10_cal = 16'b0000001110010000;
            15'd7975: log10_cal = 16'b0000001110010000;
            15'd7976: log10_cal = 16'b0000001110010000;
            15'd7977: log10_cal = 16'b0000001110010000;
            15'd7978: log10_cal = 16'b0000001110010000;
            15'd7979: log10_cal = 16'b0000001110010001;
            15'd7980: log10_cal = 16'b0000001110010001;
            15'd7981: log10_cal = 16'b0000001110010001;
            15'd7982: log10_cal = 16'b0000001110010001;
            15'd7983: log10_cal = 16'b0000001110010001;
            15'd7984: log10_cal = 16'b0000001110010001;
            15'd7985: log10_cal = 16'b0000001110010001;
            15'd7986: log10_cal = 16'b0000001110010001;
            15'd7987: log10_cal = 16'b0000001110010001;
            15'd7988: log10_cal = 16'b0000001110010001;
            15'd7989: log10_cal = 16'b0000001110010001;
            15'd7990: log10_cal = 16'b0000001110010001;
            15'd7991: log10_cal = 16'b0000001110010001;
            15'd7992: log10_cal = 16'b0000001110010001;
            15'd7993: log10_cal = 16'b0000001110010001;
            15'd7994: log10_cal = 16'b0000001110010001;
            15'd7995: log10_cal = 16'b0000001110010001;
            15'd7996: log10_cal = 16'b0000001110010001;
            15'd7997: log10_cal = 16'b0000001110010010;
            15'd7998: log10_cal = 16'b0000001110010010;
            15'd7999: log10_cal = 16'b0000001110010010;
            15'd8000: log10_cal = 16'b0000001110010010;
            15'd8001: log10_cal = 16'b0000001110010010;
            15'd8002: log10_cal = 16'b0000001110010010;
            15'd8003: log10_cal = 16'b0000001110010010;
            15'd8004: log10_cal = 16'b0000001110010010;
            15'd8005: log10_cal = 16'b0000001110010010;
            15'd8006: log10_cal = 16'b0000001110010010;
            15'd8007: log10_cal = 16'b0000001110010010;
            15'd8008: log10_cal = 16'b0000001110010010;
            15'd8009: log10_cal = 16'b0000001110010010;
            15'd8010: log10_cal = 16'b0000001110010010;
            15'd8011: log10_cal = 16'b0000001110010010;
            15'd8012: log10_cal = 16'b0000001110010010;
            15'd8013: log10_cal = 16'b0000001110010010;
            15'd8014: log10_cal = 16'b0000001110010010;
            15'd8015: log10_cal = 16'b0000001110010011;
            15'd8016: log10_cal = 16'b0000001110010011;
            15'd8017: log10_cal = 16'b0000001110010011;
            15'd8018: log10_cal = 16'b0000001110010011;
            15'd8019: log10_cal = 16'b0000001110010011;
            15'd8020: log10_cal = 16'b0000001110010011;
            15'd8021: log10_cal = 16'b0000001110010011;
            15'd8022: log10_cal = 16'b0000001110010011;
            15'd8023: log10_cal = 16'b0000001110010011;
            15'd8024: log10_cal = 16'b0000001110010011;
            15'd8025: log10_cal = 16'b0000001110010011;
            15'd8026: log10_cal = 16'b0000001110010011;
            15'd8027: log10_cal = 16'b0000001110010011;
            15'd8028: log10_cal = 16'b0000001110010011;
            15'd8029: log10_cal = 16'b0000001110010011;
            15'd8030: log10_cal = 16'b0000001110010011;
            15'd8031: log10_cal = 16'b0000001110010011;
            15'd8032: log10_cal = 16'b0000001110010011;
            15'd8033: log10_cal = 16'b0000001110010100;
            15'd8034: log10_cal = 16'b0000001110010100;
            15'd8035: log10_cal = 16'b0000001110010100;
            15'd8036: log10_cal = 16'b0000001110010100;
            15'd8037: log10_cal = 16'b0000001110010100;
            15'd8038: log10_cal = 16'b0000001110010100;
            15'd8039: log10_cal = 16'b0000001110010100;
            15'd8040: log10_cal = 16'b0000001110010100;
            15'd8041: log10_cal = 16'b0000001110010100;
            15'd8042: log10_cal = 16'b0000001110010100;
            15'd8043: log10_cal = 16'b0000001110010100;
            15'd8044: log10_cal = 16'b0000001110010100;
            15'd8045: log10_cal = 16'b0000001110010100;
            15'd8046: log10_cal = 16'b0000001110010100;
            15'd8047: log10_cal = 16'b0000001110010100;
            15'd8048: log10_cal = 16'b0000001110010100;
            15'd8049: log10_cal = 16'b0000001110010100;
            15'd8050: log10_cal = 16'b0000001110010100;
            15'd8051: log10_cal = 16'b0000001110010101;
            15'd8052: log10_cal = 16'b0000001110010101;
            15'd8053: log10_cal = 16'b0000001110010101;
            15'd8054: log10_cal = 16'b0000001110010101;
            15'd8055: log10_cal = 16'b0000001110010101;
            15'd8056: log10_cal = 16'b0000001110010101;
            15'd8057: log10_cal = 16'b0000001110010101;
            15'd8058: log10_cal = 16'b0000001110010101;
            15'd8059: log10_cal = 16'b0000001110010101;
            15'd8060: log10_cal = 16'b0000001110010101;
            15'd8061: log10_cal = 16'b0000001110010101;
            15'd8062: log10_cal = 16'b0000001110010101;
            15'd8063: log10_cal = 16'b0000001110010101;
            15'd8064: log10_cal = 16'b0000001110010101;
            15'd8065: log10_cal = 16'b0000001110010101;
            15'd8066: log10_cal = 16'b0000001110010101;
            15'd8067: log10_cal = 16'b0000001110010101;
            15'd8068: log10_cal = 16'b0000001110010101;
            15'd8069: log10_cal = 16'b0000001110010110;
            15'd8070: log10_cal = 16'b0000001110010110;
            15'd8071: log10_cal = 16'b0000001110010110;
            15'd8072: log10_cal = 16'b0000001110010110;
            15'd8073: log10_cal = 16'b0000001110010110;
            15'd8074: log10_cal = 16'b0000001110010110;
            15'd8075: log10_cal = 16'b0000001110010110;
            15'd8076: log10_cal = 16'b0000001110010110;
            15'd8077: log10_cal = 16'b0000001110010110;
            15'd8078: log10_cal = 16'b0000001110010110;
            15'd8079: log10_cal = 16'b0000001110010110;
            15'd8080: log10_cal = 16'b0000001110010110;
            15'd8081: log10_cal = 16'b0000001110010110;
            15'd8082: log10_cal = 16'b0000001110010110;
            15'd8083: log10_cal = 16'b0000001110010110;
            15'd8084: log10_cal = 16'b0000001110010110;
            15'd8085: log10_cal = 16'b0000001110010110;
            15'd8086: log10_cal = 16'b0000001110010110;
            15'd8087: log10_cal = 16'b0000001110010111;
            15'd8088: log10_cal = 16'b0000001110010111;
            15'd8089: log10_cal = 16'b0000001110010111;
            15'd8090: log10_cal = 16'b0000001110010111;
            15'd8091: log10_cal = 16'b0000001110010111;
            15'd8092: log10_cal = 16'b0000001110010111;
            15'd8093: log10_cal = 16'b0000001110010111;
            15'd8094: log10_cal = 16'b0000001110010111;
            15'd8095: log10_cal = 16'b0000001110010111;
            15'd8096: log10_cal = 16'b0000001110010111;
            15'd8097: log10_cal = 16'b0000001110010111;
            15'd8098: log10_cal = 16'b0000001110010111;
            15'd8099: log10_cal = 16'b0000001110010111;
            15'd8100: log10_cal = 16'b0000001110010111;
            15'd8101: log10_cal = 16'b0000001110010111;
            15'd8102: log10_cal = 16'b0000001110010111;
            15'd8103: log10_cal = 16'b0000001110010111;
            15'd8104: log10_cal = 16'b0000001110010111;
            15'd8105: log10_cal = 16'b0000001110011000;
            15'd8106: log10_cal = 16'b0000001110011000;
            15'd8107: log10_cal = 16'b0000001110011000;
            15'd8108: log10_cal = 16'b0000001110011000;
            15'd8109: log10_cal = 16'b0000001110011000;
            15'd8110: log10_cal = 16'b0000001110011000;
            15'd8111: log10_cal = 16'b0000001110011000;
            15'd8112: log10_cal = 16'b0000001110011000;
            15'd8113: log10_cal = 16'b0000001110011000;
            15'd8114: log10_cal = 16'b0000001110011000;
            15'd8115: log10_cal = 16'b0000001110011000;
            15'd8116: log10_cal = 16'b0000001110011000;
            15'd8117: log10_cal = 16'b0000001110011000;
            15'd8118: log10_cal = 16'b0000001110011000;
            15'd8119: log10_cal = 16'b0000001110011000;
            15'd8120: log10_cal = 16'b0000001110011000;
            15'd8121: log10_cal = 16'b0000001110011000;
            15'd8122: log10_cal = 16'b0000001110011000;
            15'd8123: log10_cal = 16'b0000001110011001;
            15'd8124: log10_cal = 16'b0000001110011001;
            15'd8125: log10_cal = 16'b0000001110011001;
            15'd8126: log10_cal = 16'b0000001110011001;
            15'd8127: log10_cal = 16'b0000001110011001;
            15'd8128: log10_cal = 16'b0000001110011001;
            15'd8129: log10_cal = 16'b0000001110011001;
            15'd8130: log10_cal = 16'b0000001110011001;
            15'd8131: log10_cal = 16'b0000001110011001;
            15'd8132: log10_cal = 16'b0000001110011001;
            15'd8133: log10_cal = 16'b0000001110011001;
            15'd8134: log10_cal = 16'b0000001110011001;
            15'd8135: log10_cal = 16'b0000001110011001;
            15'd8136: log10_cal = 16'b0000001110011001;
            15'd8137: log10_cal = 16'b0000001110011001;
            15'd8138: log10_cal = 16'b0000001110011001;
            15'd8139: log10_cal = 16'b0000001110011001;
            15'd8140: log10_cal = 16'b0000001110011001;
            15'd8141: log10_cal = 16'b0000001110011001;
            15'd8142: log10_cal = 16'b0000001110011010;
            15'd8143: log10_cal = 16'b0000001110011010;
            15'd8144: log10_cal = 16'b0000001110011010;
            15'd8145: log10_cal = 16'b0000001110011010;
            15'd8146: log10_cal = 16'b0000001110011010;
            15'd8147: log10_cal = 16'b0000001110011010;
            15'd8148: log10_cal = 16'b0000001110011010;
            15'd8149: log10_cal = 16'b0000001110011010;
            15'd8150: log10_cal = 16'b0000001110011010;
            15'd8151: log10_cal = 16'b0000001110011010;
            15'd8152: log10_cal = 16'b0000001110011010;
            15'd8153: log10_cal = 16'b0000001110011010;
            15'd8154: log10_cal = 16'b0000001110011010;
            15'd8155: log10_cal = 16'b0000001110011010;
            15'd8156: log10_cal = 16'b0000001110011010;
            15'd8157: log10_cal = 16'b0000001110011010;
            15'd8158: log10_cal = 16'b0000001110011010;
            15'd8159: log10_cal = 16'b0000001110011010;
            15'd8160: log10_cal = 16'b0000001110011011;
            15'd8161: log10_cal = 16'b0000001110011011;
            15'd8162: log10_cal = 16'b0000001110011011;
            15'd8163: log10_cal = 16'b0000001110011011;
            15'd8164: log10_cal = 16'b0000001110011011;
            15'd8165: log10_cal = 16'b0000001110011011;
            15'd8166: log10_cal = 16'b0000001110011011;
            15'd8167: log10_cal = 16'b0000001110011011;
            15'd8168: log10_cal = 16'b0000001110011011;
            15'd8169: log10_cal = 16'b0000001110011011;
            15'd8170: log10_cal = 16'b0000001110011011;
            15'd8171: log10_cal = 16'b0000001110011011;
            15'd8172: log10_cal = 16'b0000001110011011;
            15'd8173: log10_cal = 16'b0000001110011011;
            15'd8174: log10_cal = 16'b0000001110011011;
            15'd8175: log10_cal = 16'b0000001110011011;
            15'd8176: log10_cal = 16'b0000001110011011;
            15'd8177: log10_cal = 16'b0000001110011011;
            15'd8178: log10_cal = 16'b0000001110011100;
            15'd8179: log10_cal = 16'b0000001110011100;
            15'd8180: log10_cal = 16'b0000001110011100;
            15'd8181: log10_cal = 16'b0000001110011100;
            15'd8182: log10_cal = 16'b0000001110011100;
            15'd8183: log10_cal = 16'b0000001110011100;
            15'd8184: log10_cal = 16'b0000001110011100;
            15'd8185: log10_cal = 16'b0000001110011100;
            15'd8186: log10_cal = 16'b0000001110011100;
            15'd8187: log10_cal = 16'b0000001110011100;
            15'd8188: log10_cal = 16'b0000001110011100;
            15'd8189: log10_cal = 16'b0000001110011100;
            15'd8190: log10_cal = 16'b0000001110011100;
            15'd8191: log10_cal = 16'b0000001110011100;
            15'd8192: log10_cal = 16'b0000001110011100;
            15'd8193: log10_cal = 16'b0000001110011100;
            15'd8194: log10_cal = 16'b0000001110011100;
            15'd8195: log10_cal = 16'b0000001110011100;
            15'd8196: log10_cal = 16'b0000001110011100;
            15'd8197: log10_cal = 16'b0000001110011101;
            15'd8198: log10_cal = 16'b0000001110011101;
            15'd8199: log10_cal = 16'b0000001110011101;
            15'd8200: log10_cal = 16'b0000001110011101;
            15'd8201: log10_cal = 16'b0000001110011101;
            15'd8202: log10_cal = 16'b0000001110011101;
            15'd8203: log10_cal = 16'b0000001110011101;
            15'd8204: log10_cal = 16'b0000001110011101;
            15'd8205: log10_cal = 16'b0000001110011101;
            15'd8206: log10_cal = 16'b0000001110011101;
            15'd8207: log10_cal = 16'b0000001110011101;
            15'd8208: log10_cal = 16'b0000001110011101;
            15'd8209: log10_cal = 16'b0000001110011101;
            15'd8210: log10_cal = 16'b0000001110011101;
            15'd8211: log10_cal = 16'b0000001110011101;
            15'd8212: log10_cal = 16'b0000001110011101;
            15'd8213: log10_cal = 16'b0000001110011101;
            15'd8214: log10_cal = 16'b0000001110011101;
            15'd8215: log10_cal = 16'b0000001110011110;
            15'd8216: log10_cal = 16'b0000001110011110;
            15'd8217: log10_cal = 16'b0000001110011110;
            15'd8218: log10_cal = 16'b0000001110011110;
            15'd8219: log10_cal = 16'b0000001110011110;
            15'd8220: log10_cal = 16'b0000001110011110;
            15'd8221: log10_cal = 16'b0000001110011110;
            15'd8222: log10_cal = 16'b0000001110011110;
            15'd8223: log10_cal = 16'b0000001110011110;
            15'd8224: log10_cal = 16'b0000001110011110;
            15'd8225: log10_cal = 16'b0000001110011110;
            15'd8226: log10_cal = 16'b0000001110011110;
            15'd8227: log10_cal = 16'b0000001110011110;
            15'd8228: log10_cal = 16'b0000001110011110;
            15'd8229: log10_cal = 16'b0000001110011110;
            15'd8230: log10_cal = 16'b0000001110011110;
            15'd8231: log10_cal = 16'b0000001110011110;
            15'd8232: log10_cal = 16'b0000001110011110;
            15'd8233: log10_cal = 16'b0000001110011110;
            15'd8234: log10_cal = 16'b0000001110011111;
            15'd8235: log10_cal = 16'b0000001110011111;
            15'd8236: log10_cal = 16'b0000001110011111;
            15'd8237: log10_cal = 16'b0000001110011111;
            15'd8238: log10_cal = 16'b0000001110011111;
            15'd8239: log10_cal = 16'b0000001110011111;
            15'd8240: log10_cal = 16'b0000001110011111;
            15'd8241: log10_cal = 16'b0000001110011111;
            15'd8242: log10_cal = 16'b0000001110011111;
            15'd8243: log10_cal = 16'b0000001110011111;
            15'd8244: log10_cal = 16'b0000001110011111;
            15'd8245: log10_cal = 16'b0000001110011111;
            15'd8246: log10_cal = 16'b0000001110011111;
            15'd8247: log10_cal = 16'b0000001110011111;
            15'd8248: log10_cal = 16'b0000001110011111;
            15'd8249: log10_cal = 16'b0000001110011111;
            15'd8250: log10_cal = 16'b0000001110011111;
            15'd8251: log10_cal = 16'b0000001110011111;
            15'd8252: log10_cal = 16'b0000001110100000;
            15'd8253: log10_cal = 16'b0000001110100000;
            15'd8254: log10_cal = 16'b0000001110100000;
            15'd8255: log10_cal = 16'b0000001110100000;
            15'd8256: log10_cal = 16'b0000001110100000;
            15'd8257: log10_cal = 16'b0000001110100000;
            15'd8258: log10_cal = 16'b0000001110100000;
            15'd8259: log10_cal = 16'b0000001110100000;
            15'd8260: log10_cal = 16'b0000001110100000;
            15'd8261: log10_cal = 16'b0000001110100000;
            15'd8262: log10_cal = 16'b0000001110100000;
            15'd8263: log10_cal = 16'b0000001110100000;
            15'd8264: log10_cal = 16'b0000001110100000;
            15'd8265: log10_cal = 16'b0000001110100000;
            15'd8266: log10_cal = 16'b0000001110100000;
            15'd8267: log10_cal = 16'b0000001110100000;
            15'd8268: log10_cal = 16'b0000001110100000;
            15'd8269: log10_cal = 16'b0000001110100000;
            15'd8270: log10_cal = 16'b0000001110100000;
            15'd8271: log10_cal = 16'b0000001110100001;
            15'd8272: log10_cal = 16'b0000001110100001;
            15'd8273: log10_cal = 16'b0000001110100001;
            15'd8274: log10_cal = 16'b0000001110100001;
            15'd8275: log10_cal = 16'b0000001110100001;
            15'd8276: log10_cal = 16'b0000001110100001;
            15'd8277: log10_cal = 16'b0000001110100001;
            15'd8278: log10_cal = 16'b0000001110100001;
            15'd8279: log10_cal = 16'b0000001110100001;
            15'd8280: log10_cal = 16'b0000001110100001;
            15'd8281: log10_cal = 16'b0000001110100001;
            15'd8282: log10_cal = 16'b0000001110100001;
            15'd8283: log10_cal = 16'b0000001110100001;
            15'd8284: log10_cal = 16'b0000001110100001;
            15'd8285: log10_cal = 16'b0000001110100001;
            15'd8286: log10_cal = 16'b0000001110100001;
            15'd8287: log10_cal = 16'b0000001110100001;
            15'd8288: log10_cal = 16'b0000001110100001;
            15'd8289: log10_cal = 16'b0000001110100001;
            15'd8290: log10_cal = 16'b0000001110100010;
            15'd8291: log10_cal = 16'b0000001110100010;
            15'd8292: log10_cal = 16'b0000001110100010;
            15'd8293: log10_cal = 16'b0000001110100010;
            15'd8294: log10_cal = 16'b0000001110100010;
            15'd8295: log10_cal = 16'b0000001110100010;
            15'd8296: log10_cal = 16'b0000001110100010;
            15'd8297: log10_cal = 16'b0000001110100010;
            15'd8298: log10_cal = 16'b0000001110100010;
            15'd8299: log10_cal = 16'b0000001110100010;
            15'd8300: log10_cal = 16'b0000001110100010;
            15'd8301: log10_cal = 16'b0000001110100010;
            15'd8302: log10_cal = 16'b0000001110100010;
            15'd8303: log10_cal = 16'b0000001110100010;
            15'd8304: log10_cal = 16'b0000001110100010;
            15'd8305: log10_cal = 16'b0000001110100010;
            15'd8306: log10_cal = 16'b0000001110100010;
            15'd8307: log10_cal = 16'b0000001110100010;
            15'd8308: log10_cal = 16'b0000001110100011;
            15'd8309: log10_cal = 16'b0000001110100011;
            15'd8310: log10_cal = 16'b0000001110100011;
            15'd8311: log10_cal = 16'b0000001110100011;
            15'd8312: log10_cal = 16'b0000001110100011;
            15'd8313: log10_cal = 16'b0000001110100011;
            15'd8314: log10_cal = 16'b0000001110100011;
            15'd8315: log10_cal = 16'b0000001110100011;
            15'd8316: log10_cal = 16'b0000001110100011;
            15'd8317: log10_cal = 16'b0000001110100011;
            15'd8318: log10_cal = 16'b0000001110100011;
            15'd8319: log10_cal = 16'b0000001110100011;
            15'd8320: log10_cal = 16'b0000001110100011;
            15'd8321: log10_cal = 16'b0000001110100011;
            15'd8322: log10_cal = 16'b0000001110100011;
            15'd8323: log10_cal = 16'b0000001110100011;
            15'd8324: log10_cal = 16'b0000001110100011;
            15'd8325: log10_cal = 16'b0000001110100011;
            15'd8326: log10_cal = 16'b0000001110100011;
            15'd8327: log10_cal = 16'b0000001110100100;
            15'd8328: log10_cal = 16'b0000001110100100;
            15'd8329: log10_cal = 16'b0000001110100100;
            15'd8330: log10_cal = 16'b0000001110100100;
            15'd8331: log10_cal = 16'b0000001110100100;
            15'd8332: log10_cal = 16'b0000001110100100;
            15'd8333: log10_cal = 16'b0000001110100100;
            15'd8334: log10_cal = 16'b0000001110100100;
            15'd8335: log10_cal = 16'b0000001110100100;
            15'd8336: log10_cal = 16'b0000001110100100;
            15'd8337: log10_cal = 16'b0000001110100100;
            15'd8338: log10_cal = 16'b0000001110100100;
            15'd8339: log10_cal = 16'b0000001110100100;
            15'd8340: log10_cal = 16'b0000001110100100;
            15'd8341: log10_cal = 16'b0000001110100100;
            15'd8342: log10_cal = 16'b0000001110100100;
            15'd8343: log10_cal = 16'b0000001110100100;
            15'd8344: log10_cal = 16'b0000001110100100;
            15'd8345: log10_cal = 16'b0000001110100100;
            15'd8346: log10_cal = 16'b0000001110100101;
            15'd8347: log10_cal = 16'b0000001110100101;
            15'd8348: log10_cal = 16'b0000001110100101;
            15'd8349: log10_cal = 16'b0000001110100101;
            15'd8350: log10_cal = 16'b0000001110100101;
            15'd8351: log10_cal = 16'b0000001110100101;
            15'd8352: log10_cal = 16'b0000001110100101;
            15'd8353: log10_cal = 16'b0000001110100101;
            15'd8354: log10_cal = 16'b0000001110100101;
            15'd8355: log10_cal = 16'b0000001110100101;
            15'd8356: log10_cal = 16'b0000001110100101;
            15'd8357: log10_cal = 16'b0000001110100101;
            15'd8358: log10_cal = 16'b0000001110100101;
            15'd8359: log10_cal = 16'b0000001110100101;
            15'd8360: log10_cal = 16'b0000001110100101;
            15'd8361: log10_cal = 16'b0000001110100101;
            15'd8362: log10_cal = 16'b0000001110100101;
            15'd8363: log10_cal = 16'b0000001110100101;
            15'd8364: log10_cal = 16'b0000001110100110;
            15'd8365: log10_cal = 16'b0000001110100110;
            15'd8366: log10_cal = 16'b0000001110100110;
            15'd8367: log10_cal = 16'b0000001110100110;
            15'd8368: log10_cal = 16'b0000001110100110;
            15'd8369: log10_cal = 16'b0000001110100110;
            15'd8370: log10_cal = 16'b0000001110100110;
            15'd8371: log10_cal = 16'b0000001110100110;
            15'd8372: log10_cal = 16'b0000001110100110;
            15'd8373: log10_cal = 16'b0000001110100110;
            15'd8374: log10_cal = 16'b0000001110100110;
            15'd8375: log10_cal = 16'b0000001110100110;
            15'd8376: log10_cal = 16'b0000001110100110;
            15'd8377: log10_cal = 16'b0000001110100110;
            15'd8378: log10_cal = 16'b0000001110100110;
            15'd8379: log10_cal = 16'b0000001110100110;
            15'd8380: log10_cal = 16'b0000001110100110;
            15'd8381: log10_cal = 16'b0000001110100110;
            15'd8382: log10_cal = 16'b0000001110100110;
            15'd8383: log10_cal = 16'b0000001110100111;
            15'd8384: log10_cal = 16'b0000001110100111;
            15'd8385: log10_cal = 16'b0000001110100111;
            15'd8386: log10_cal = 16'b0000001110100111;
            15'd8387: log10_cal = 16'b0000001110100111;
            15'd8388: log10_cal = 16'b0000001110100111;
            15'd8389: log10_cal = 16'b0000001110100111;
            15'd8390: log10_cal = 16'b0000001110100111;
            15'd8391: log10_cal = 16'b0000001110100111;
            15'd8392: log10_cal = 16'b0000001110100111;
            15'd8393: log10_cal = 16'b0000001110100111;
            15'd8394: log10_cal = 16'b0000001110100111;
            15'd8395: log10_cal = 16'b0000001110100111;
            15'd8396: log10_cal = 16'b0000001110100111;
            15'd8397: log10_cal = 16'b0000001110100111;
            15'd8398: log10_cal = 16'b0000001110100111;
            15'd8399: log10_cal = 16'b0000001110100111;
            15'd8400: log10_cal = 16'b0000001110100111;
            15'd8401: log10_cal = 16'b0000001110100111;
            15'd8402: log10_cal = 16'b0000001110101000;
            15'd8403: log10_cal = 16'b0000001110101000;
            15'd8404: log10_cal = 16'b0000001110101000;
            15'd8405: log10_cal = 16'b0000001110101000;
            15'd8406: log10_cal = 16'b0000001110101000;
            15'd8407: log10_cal = 16'b0000001110101000;
            15'd8408: log10_cal = 16'b0000001110101000;
            15'd8409: log10_cal = 16'b0000001110101000;
            15'd8410: log10_cal = 16'b0000001110101000;
            15'd8411: log10_cal = 16'b0000001110101000;
            15'd8412: log10_cal = 16'b0000001110101000;
            15'd8413: log10_cal = 16'b0000001110101000;
            15'd8414: log10_cal = 16'b0000001110101000;
            15'd8415: log10_cal = 16'b0000001110101000;
            15'd8416: log10_cal = 16'b0000001110101000;
            15'd8417: log10_cal = 16'b0000001110101000;
            15'd8418: log10_cal = 16'b0000001110101000;
            15'd8419: log10_cal = 16'b0000001110101000;
            15'd8420: log10_cal = 16'b0000001110101000;
            15'd8421: log10_cal = 16'b0000001110101001;
            15'd8422: log10_cal = 16'b0000001110101001;
            15'd8423: log10_cal = 16'b0000001110101001;
            15'd8424: log10_cal = 16'b0000001110101001;
            15'd8425: log10_cal = 16'b0000001110101001;
            15'd8426: log10_cal = 16'b0000001110101001;
            15'd8427: log10_cal = 16'b0000001110101001;
            15'd8428: log10_cal = 16'b0000001110101001;
            15'd8429: log10_cal = 16'b0000001110101001;
            15'd8430: log10_cal = 16'b0000001110101001;
            15'd8431: log10_cal = 16'b0000001110101001;
            15'd8432: log10_cal = 16'b0000001110101001;
            15'd8433: log10_cal = 16'b0000001110101001;
            15'd8434: log10_cal = 16'b0000001110101001;
            15'd8435: log10_cal = 16'b0000001110101001;
            15'd8436: log10_cal = 16'b0000001110101001;
            15'd8437: log10_cal = 16'b0000001110101001;
            15'd8438: log10_cal = 16'b0000001110101001;
            15'd8439: log10_cal = 16'b0000001110101001;
            15'd8440: log10_cal = 16'b0000001110101010;
            15'd8441: log10_cal = 16'b0000001110101010;
            15'd8442: log10_cal = 16'b0000001110101010;
            15'd8443: log10_cal = 16'b0000001110101010;
            15'd8444: log10_cal = 16'b0000001110101010;
            15'd8445: log10_cal = 16'b0000001110101010;
            15'd8446: log10_cal = 16'b0000001110101010;
            15'd8447: log10_cal = 16'b0000001110101010;
            15'd8448: log10_cal = 16'b0000001110101010;
            15'd8449: log10_cal = 16'b0000001110101010;
            15'd8450: log10_cal = 16'b0000001110101010;
            15'd8451: log10_cal = 16'b0000001110101010;
            15'd8452: log10_cal = 16'b0000001110101010;
            15'd8453: log10_cal = 16'b0000001110101010;
            15'd8454: log10_cal = 16'b0000001110101010;
            15'd8455: log10_cal = 16'b0000001110101010;
            15'd8456: log10_cal = 16'b0000001110101010;
            15'd8457: log10_cal = 16'b0000001110101010;
            15'd8458: log10_cal = 16'b0000001110101010;
            15'd8459: log10_cal = 16'b0000001110101011;
            15'd8460: log10_cal = 16'b0000001110101011;
            15'd8461: log10_cal = 16'b0000001110101011;
            15'd8462: log10_cal = 16'b0000001110101011;
            15'd8463: log10_cal = 16'b0000001110101011;
            15'd8464: log10_cal = 16'b0000001110101011;
            15'd8465: log10_cal = 16'b0000001110101011;
            15'd8466: log10_cal = 16'b0000001110101011;
            15'd8467: log10_cal = 16'b0000001110101011;
            15'd8468: log10_cal = 16'b0000001110101011;
            15'd8469: log10_cal = 16'b0000001110101011;
            15'd8470: log10_cal = 16'b0000001110101011;
            15'd8471: log10_cal = 16'b0000001110101011;
            15'd8472: log10_cal = 16'b0000001110101011;
            15'd8473: log10_cal = 16'b0000001110101011;
            15'd8474: log10_cal = 16'b0000001110101011;
            15'd8475: log10_cal = 16'b0000001110101011;
            15'd8476: log10_cal = 16'b0000001110101011;
            15'd8477: log10_cal = 16'b0000001110101011;
            15'd8478: log10_cal = 16'b0000001110101100;
            15'd8479: log10_cal = 16'b0000001110101100;
            15'd8480: log10_cal = 16'b0000001110101100;
            15'd8481: log10_cal = 16'b0000001110101100;
            15'd8482: log10_cal = 16'b0000001110101100;
            15'd8483: log10_cal = 16'b0000001110101100;
            15'd8484: log10_cal = 16'b0000001110101100;
            15'd8485: log10_cal = 16'b0000001110101100;
            15'd8486: log10_cal = 16'b0000001110101100;
            15'd8487: log10_cal = 16'b0000001110101100;
            15'd8488: log10_cal = 16'b0000001110101100;
            15'd8489: log10_cal = 16'b0000001110101100;
            15'd8490: log10_cal = 16'b0000001110101100;
            15'd8491: log10_cal = 16'b0000001110101100;
            15'd8492: log10_cal = 16'b0000001110101100;
            15'd8493: log10_cal = 16'b0000001110101100;
            15'd8494: log10_cal = 16'b0000001110101100;
            15'd8495: log10_cal = 16'b0000001110101100;
            15'd8496: log10_cal = 16'b0000001110101100;
            15'd8497: log10_cal = 16'b0000001110101101;
            15'd8498: log10_cal = 16'b0000001110101101;
            15'd8499: log10_cal = 16'b0000001110101101;
            15'd8500: log10_cal = 16'b0000001110101101;
            15'd8501: log10_cal = 16'b0000001110101101;
            15'd8502: log10_cal = 16'b0000001110101101;
            15'd8503: log10_cal = 16'b0000001110101101;
            15'd8504: log10_cal = 16'b0000001110101101;
            15'd8505: log10_cal = 16'b0000001110101101;
            15'd8506: log10_cal = 16'b0000001110101101;
            15'd8507: log10_cal = 16'b0000001110101101;
            15'd8508: log10_cal = 16'b0000001110101101;
            15'd8509: log10_cal = 16'b0000001110101101;
            15'd8510: log10_cal = 16'b0000001110101101;
            15'd8511: log10_cal = 16'b0000001110101101;
            15'd8512: log10_cal = 16'b0000001110101101;
            15'd8513: log10_cal = 16'b0000001110101101;
            15'd8514: log10_cal = 16'b0000001110101101;
            15'd8515: log10_cal = 16'b0000001110101101;
            15'd8516: log10_cal = 16'b0000001110101110;
            15'd8517: log10_cal = 16'b0000001110101110;
            15'd8518: log10_cal = 16'b0000001110101110;
            15'd8519: log10_cal = 16'b0000001110101110;
            15'd8520: log10_cal = 16'b0000001110101110;
            15'd8521: log10_cal = 16'b0000001110101110;
            15'd8522: log10_cal = 16'b0000001110101110;
            15'd8523: log10_cal = 16'b0000001110101110;
            15'd8524: log10_cal = 16'b0000001110101110;
            15'd8525: log10_cal = 16'b0000001110101110;
            15'd8526: log10_cal = 16'b0000001110101110;
            15'd8527: log10_cal = 16'b0000001110101110;
            15'd8528: log10_cal = 16'b0000001110101110;
            15'd8529: log10_cal = 16'b0000001110101110;
            15'd8530: log10_cal = 16'b0000001110101110;
            15'd8531: log10_cal = 16'b0000001110101110;
            15'd8532: log10_cal = 16'b0000001110101110;
            15'd8533: log10_cal = 16'b0000001110101110;
            15'd8534: log10_cal = 16'b0000001110101110;
            15'd8535: log10_cal = 16'b0000001110101111;
            15'd8536: log10_cal = 16'b0000001110101111;
            15'd8537: log10_cal = 16'b0000001110101111;
            15'd8538: log10_cal = 16'b0000001110101111;
            15'd8539: log10_cal = 16'b0000001110101111;
            15'd8540: log10_cal = 16'b0000001110101111;
            15'd8541: log10_cal = 16'b0000001110101111;
            15'd8542: log10_cal = 16'b0000001110101111;
            15'd8543: log10_cal = 16'b0000001110101111;
            15'd8544: log10_cal = 16'b0000001110101111;
            15'd8545: log10_cal = 16'b0000001110101111;
            15'd8546: log10_cal = 16'b0000001110101111;
            15'd8547: log10_cal = 16'b0000001110101111;
            15'd8548: log10_cal = 16'b0000001110101111;
            15'd8549: log10_cal = 16'b0000001110101111;
            15'd8550: log10_cal = 16'b0000001110101111;
            15'd8551: log10_cal = 16'b0000001110101111;
            15'd8552: log10_cal = 16'b0000001110101111;
            15'd8553: log10_cal = 16'b0000001110101111;
            15'd8554: log10_cal = 16'b0000001110101111;
            15'd8555: log10_cal = 16'b0000001110110000;
            15'd8556: log10_cal = 16'b0000001110110000;
            15'd8557: log10_cal = 16'b0000001110110000;
            15'd8558: log10_cal = 16'b0000001110110000;
            15'd8559: log10_cal = 16'b0000001110110000;
            15'd8560: log10_cal = 16'b0000001110110000;
            15'd8561: log10_cal = 16'b0000001110110000;
            15'd8562: log10_cal = 16'b0000001110110000;
            15'd8563: log10_cal = 16'b0000001110110000;
            15'd8564: log10_cal = 16'b0000001110110000;
            15'd8565: log10_cal = 16'b0000001110110000;
            15'd8566: log10_cal = 16'b0000001110110000;
            15'd8567: log10_cal = 16'b0000001110110000;
            15'd8568: log10_cal = 16'b0000001110110000;
            15'd8569: log10_cal = 16'b0000001110110000;
            15'd8570: log10_cal = 16'b0000001110110000;
            15'd8571: log10_cal = 16'b0000001110110000;
            15'd8572: log10_cal = 16'b0000001110110000;
            15'd8573: log10_cal = 16'b0000001110110000;
            15'd8574: log10_cal = 16'b0000001110110001;
            15'd8575: log10_cal = 16'b0000001110110001;
            15'd8576: log10_cal = 16'b0000001110110001;
            15'd8577: log10_cal = 16'b0000001110110001;
            15'd8578: log10_cal = 16'b0000001110110001;
            15'd8579: log10_cal = 16'b0000001110110001;
            15'd8580: log10_cal = 16'b0000001110110001;
            15'd8581: log10_cal = 16'b0000001110110001;
            15'd8582: log10_cal = 16'b0000001110110001;
            15'd8583: log10_cal = 16'b0000001110110001;
            15'd8584: log10_cal = 16'b0000001110110001;
            15'd8585: log10_cal = 16'b0000001110110001;
            15'd8586: log10_cal = 16'b0000001110110001;
            15'd8587: log10_cal = 16'b0000001110110001;
            15'd8588: log10_cal = 16'b0000001110110001;
            15'd8589: log10_cal = 16'b0000001110110001;
            15'd8590: log10_cal = 16'b0000001110110001;
            15'd8591: log10_cal = 16'b0000001110110001;
            15'd8592: log10_cal = 16'b0000001110110001;
            15'd8593: log10_cal = 16'b0000001110110010;
            15'd8594: log10_cal = 16'b0000001110110010;
            15'd8595: log10_cal = 16'b0000001110110010;
            15'd8596: log10_cal = 16'b0000001110110010;
            15'd8597: log10_cal = 16'b0000001110110010;
            15'd8598: log10_cal = 16'b0000001110110010;
            15'd8599: log10_cal = 16'b0000001110110010;
            15'd8600: log10_cal = 16'b0000001110110010;
            15'd8601: log10_cal = 16'b0000001110110010;
            15'd8602: log10_cal = 16'b0000001110110010;
            15'd8603: log10_cal = 16'b0000001110110010;
            15'd8604: log10_cal = 16'b0000001110110010;
            15'd8605: log10_cal = 16'b0000001110110010;
            15'd8606: log10_cal = 16'b0000001110110010;
            15'd8607: log10_cal = 16'b0000001110110010;
            15'd8608: log10_cal = 16'b0000001110110010;
            15'd8609: log10_cal = 16'b0000001110110010;
            15'd8610: log10_cal = 16'b0000001110110010;
            15'd8611: log10_cal = 16'b0000001110110010;
            15'd8612: log10_cal = 16'b0000001110110010;
            15'd8613: log10_cal = 16'b0000001110110011;
            15'd8614: log10_cal = 16'b0000001110110011;
            15'd8615: log10_cal = 16'b0000001110110011;
            15'd8616: log10_cal = 16'b0000001110110011;
            15'd8617: log10_cal = 16'b0000001110110011;
            15'd8618: log10_cal = 16'b0000001110110011;
            15'd8619: log10_cal = 16'b0000001110110011;
            15'd8620: log10_cal = 16'b0000001110110011;
            15'd8621: log10_cal = 16'b0000001110110011;
            15'd8622: log10_cal = 16'b0000001110110011;
            15'd8623: log10_cal = 16'b0000001110110011;
            15'd8624: log10_cal = 16'b0000001110110011;
            15'd8625: log10_cal = 16'b0000001110110011;
            15'd8626: log10_cal = 16'b0000001110110011;
            15'd8627: log10_cal = 16'b0000001110110011;
            15'd8628: log10_cal = 16'b0000001110110011;
            15'd8629: log10_cal = 16'b0000001110110011;
            15'd8630: log10_cal = 16'b0000001110110011;
            15'd8631: log10_cal = 16'b0000001110110011;
            15'd8632: log10_cal = 16'b0000001110110100;
            15'd8633: log10_cal = 16'b0000001110110100;
            15'd8634: log10_cal = 16'b0000001110110100;
            15'd8635: log10_cal = 16'b0000001110110100;
            15'd8636: log10_cal = 16'b0000001110110100;
            15'd8637: log10_cal = 16'b0000001110110100;
            15'd8638: log10_cal = 16'b0000001110110100;
            15'd8639: log10_cal = 16'b0000001110110100;
            15'd8640: log10_cal = 16'b0000001110110100;
            15'd8641: log10_cal = 16'b0000001110110100;
            15'd8642: log10_cal = 16'b0000001110110100;
            15'd8643: log10_cal = 16'b0000001110110100;
            15'd8644: log10_cal = 16'b0000001110110100;
            15'd8645: log10_cal = 16'b0000001110110100;
            15'd8646: log10_cal = 16'b0000001110110100;
            15'd8647: log10_cal = 16'b0000001110110100;
            15'd8648: log10_cal = 16'b0000001110110100;
            15'd8649: log10_cal = 16'b0000001110110100;
            15'd8650: log10_cal = 16'b0000001110110100;
            15'd8651: log10_cal = 16'b0000001110110101;
            15'd8652: log10_cal = 16'b0000001110110101;
            15'd8653: log10_cal = 16'b0000001110110101;
            15'd8654: log10_cal = 16'b0000001110110101;
            15'd8655: log10_cal = 16'b0000001110110101;
            15'd8656: log10_cal = 16'b0000001110110101;
            15'd8657: log10_cal = 16'b0000001110110101;
            15'd8658: log10_cal = 16'b0000001110110101;
            15'd8659: log10_cal = 16'b0000001110110101;
            15'd8660: log10_cal = 16'b0000001110110101;
            15'd8661: log10_cal = 16'b0000001110110101;
            15'd8662: log10_cal = 16'b0000001110110101;
            15'd8663: log10_cal = 16'b0000001110110101;
            15'd8664: log10_cal = 16'b0000001110110101;
            15'd8665: log10_cal = 16'b0000001110110101;
            15'd8666: log10_cal = 16'b0000001110110101;
            15'd8667: log10_cal = 16'b0000001110110101;
            15'd8668: log10_cal = 16'b0000001110110101;
            15'd8669: log10_cal = 16'b0000001110110101;
            15'd8670: log10_cal = 16'b0000001110110101;
            15'd8671: log10_cal = 16'b0000001110110110;
            15'd8672: log10_cal = 16'b0000001110110110;
            15'd8673: log10_cal = 16'b0000001110110110;
            15'd8674: log10_cal = 16'b0000001110110110;
            15'd8675: log10_cal = 16'b0000001110110110;
            15'd8676: log10_cal = 16'b0000001110110110;
            15'd8677: log10_cal = 16'b0000001110110110;
            15'd8678: log10_cal = 16'b0000001110110110;
            15'd8679: log10_cal = 16'b0000001110110110;
            15'd8680: log10_cal = 16'b0000001110110110;
            15'd8681: log10_cal = 16'b0000001110110110;
            15'd8682: log10_cal = 16'b0000001110110110;
            15'd8683: log10_cal = 16'b0000001110110110;
            15'd8684: log10_cal = 16'b0000001110110110;
            15'd8685: log10_cal = 16'b0000001110110110;
            15'd8686: log10_cal = 16'b0000001110110110;
            15'd8687: log10_cal = 16'b0000001110110110;
            15'd8688: log10_cal = 16'b0000001110110110;
            15'd8689: log10_cal = 16'b0000001110110110;
            15'd8690: log10_cal = 16'b0000001110110111;
            15'd8691: log10_cal = 16'b0000001110110111;
            15'd8692: log10_cal = 16'b0000001110110111;
            15'd8693: log10_cal = 16'b0000001110110111;
            15'd8694: log10_cal = 16'b0000001110110111;
            15'd8695: log10_cal = 16'b0000001110110111;
            15'd8696: log10_cal = 16'b0000001110110111;
            15'd8697: log10_cal = 16'b0000001110110111;
            15'd8698: log10_cal = 16'b0000001110110111;
            15'd8699: log10_cal = 16'b0000001110110111;
            15'd8700: log10_cal = 16'b0000001110110111;
            15'd8701: log10_cal = 16'b0000001110110111;
            15'd8702: log10_cal = 16'b0000001110110111;
            15'd8703: log10_cal = 16'b0000001110110111;
            15'd8704: log10_cal = 16'b0000001110110111;
            15'd8705: log10_cal = 16'b0000001110110111;
            15'd8706: log10_cal = 16'b0000001110110111;
            15'd8707: log10_cal = 16'b0000001110110111;
            15'd8708: log10_cal = 16'b0000001110110111;
            15'd8709: log10_cal = 16'b0000001110110111;
            15'd8710: log10_cal = 16'b0000001110111000;
            15'd8711: log10_cal = 16'b0000001110111000;
            15'd8712: log10_cal = 16'b0000001110111000;
            15'd8713: log10_cal = 16'b0000001110111000;
            15'd8714: log10_cal = 16'b0000001110111000;
            15'd8715: log10_cal = 16'b0000001110111000;
            15'd8716: log10_cal = 16'b0000001110111000;
            15'd8717: log10_cal = 16'b0000001110111000;
            15'd8718: log10_cal = 16'b0000001110111000;
            15'd8719: log10_cal = 16'b0000001110111000;
            15'd8720: log10_cal = 16'b0000001110111000;
            15'd8721: log10_cal = 16'b0000001110111000;
            15'd8722: log10_cal = 16'b0000001110111000;
            15'd8723: log10_cal = 16'b0000001110111000;
            15'd8724: log10_cal = 16'b0000001110111000;
            15'd8725: log10_cal = 16'b0000001110111000;
            15'd8726: log10_cal = 16'b0000001110111000;
            15'd8727: log10_cal = 16'b0000001110111000;
            15'd8728: log10_cal = 16'b0000001110111000;
            15'd8729: log10_cal = 16'b0000001110111001;
            15'd8730: log10_cal = 16'b0000001110111001;
            15'd8731: log10_cal = 16'b0000001110111001;
            15'd8732: log10_cal = 16'b0000001110111001;
            15'd8733: log10_cal = 16'b0000001110111001;
            15'd8734: log10_cal = 16'b0000001110111001;
            15'd8735: log10_cal = 16'b0000001110111001;
            15'd8736: log10_cal = 16'b0000001110111001;
            15'd8737: log10_cal = 16'b0000001110111001;
            15'd8738: log10_cal = 16'b0000001110111001;
            15'd8739: log10_cal = 16'b0000001110111001;
            15'd8740: log10_cal = 16'b0000001110111001;
            15'd8741: log10_cal = 16'b0000001110111001;
            15'd8742: log10_cal = 16'b0000001110111001;
            15'd8743: log10_cal = 16'b0000001110111001;
            15'd8744: log10_cal = 16'b0000001110111001;
            15'd8745: log10_cal = 16'b0000001110111001;
            15'd8746: log10_cal = 16'b0000001110111001;
            15'd8747: log10_cal = 16'b0000001110111001;
            15'd8748: log10_cal = 16'b0000001110111001;
            15'd8749: log10_cal = 16'b0000001110111010;
            15'd8750: log10_cal = 16'b0000001110111010;
            15'd8751: log10_cal = 16'b0000001110111010;
            15'd8752: log10_cal = 16'b0000001110111010;
            15'd8753: log10_cal = 16'b0000001110111010;
            15'd8754: log10_cal = 16'b0000001110111010;
            15'd8755: log10_cal = 16'b0000001110111010;
            15'd8756: log10_cal = 16'b0000001110111010;
            15'd8757: log10_cal = 16'b0000001110111010;
            15'd8758: log10_cal = 16'b0000001110111010;
            15'd8759: log10_cal = 16'b0000001110111010;
            15'd8760: log10_cal = 16'b0000001110111010;
            15'd8761: log10_cal = 16'b0000001110111010;
            15'd8762: log10_cal = 16'b0000001110111010;
            15'd8763: log10_cal = 16'b0000001110111010;
            15'd8764: log10_cal = 16'b0000001110111010;
            15'd8765: log10_cal = 16'b0000001110111010;
            15'd8766: log10_cal = 16'b0000001110111010;
            15'd8767: log10_cal = 16'b0000001110111010;
            15'd8768: log10_cal = 16'b0000001110111010;
            15'd8769: log10_cal = 16'b0000001110111011;
            15'd8770: log10_cal = 16'b0000001110111011;
            15'd8771: log10_cal = 16'b0000001110111011;
            15'd8772: log10_cal = 16'b0000001110111011;
            15'd8773: log10_cal = 16'b0000001110111011;
            15'd8774: log10_cal = 16'b0000001110111011;
            15'd8775: log10_cal = 16'b0000001110111011;
            15'd8776: log10_cal = 16'b0000001110111011;
            15'd8777: log10_cal = 16'b0000001110111011;
            15'd8778: log10_cal = 16'b0000001110111011;
            15'd8779: log10_cal = 16'b0000001110111011;
            15'd8780: log10_cal = 16'b0000001110111011;
            15'd8781: log10_cal = 16'b0000001110111011;
            15'd8782: log10_cal = 16'b0000001110111011;
            15'd8783: log10_cal = 16'b0000001110111011;
            15'd8784: log10_cal = 16'b0000001110111011;
            15'd8785: log10_cal = 16'b0000001110111011;
            15'd8786: log10_cal = 16'b0000001110111011;
            15'd8787: log10_cal = 16'b0000001110111011;
            15'd8788: log10_cal = 16'b0000001110111011;
            15'd8789: log10_cal = 16'b0000001110111100;
            15'd8790: log10_cal = 16'b0000001110111100;
            15'd8791: log10_cal = 16'b0000001110111100;
            15'd8792: log10_cal = 16'b0000001110111100;
            15'd8793: log10_cal = 16'b0000001110111100;
            15'd8794: log10_cal = 16'b0000001110111100;
            15'd8795: log10_cal = 16'b0000001110111100;
            15'd8796: log10_cal = 16'b0000001110111100;
            15'd8797: log10_cal = 16'b0000001110111100;
            15'd8798: log10_cal = 16'b0000001110111100;
            15'd8799: log10_cal = 16'b0000001110111100;
            15'd8800: log10_cal = 16'b0000001110111100;
            15'd8801: log10_cal = 16'b0000001110111100;
            15'd8802: log10_cal = 16'b0000001110111100;
            15'd8803: log10_cal = 16'b0000001110111100;
            15'd8804: log10_cal = 16'b0000001110111100;
            15'd8805: log10_cal = 16'b0000001110111100;
            15'd8806: log10_cal = 16'b0000001110111100;
            15'd8807: log10_cal = 16'b0000001110111100;
            15'd8808: log10_cal = 16'b0000001110111101;
            15'd8809: log10_cal = 16'b0000001110111101;
            15'd8810: log10_cal = 16'b0000001110111101;
            15'd8811: log10_cal = 16'b0000001110111101;
            15'd8812: log10_cal = 16'b0000001110111101;
            15'd8813: log10_cal = 16'b0000001110111101;
            15'd8814: log10_cal = 16'b0000001110111101;
            15'd8815: log10_cal = 16'b0000001110111101;
            15'd8816: log10_cal = 16'b0000001110111101;
            15'd8817: log10_cal = 16'b0000001110111101;
            15'd8818: log10_cal = 16'b0000001110111101;
            15'd8819: log10_cal = 16'b0000001110111101;
            15'd8820: log10_cal = 16'b0000001110111101;
            15'd8821: log10_cal = 16'b0000001110111101;
            15'd8822: log10_cal = 16'b0000001110111101;
            15'd8823: log10_cal = 16'b0000001110111101;
            15'd8824: log10_cal = 16'b0000001110111101;
            15'd8825: log10_cal = 16'b0000001110111101;
            15'd8826: log10_cal = 16'b0000001110111101;
            15'd8827: log10_cal = 16'b0000001110111101;
            15'd8828: log10_cal = 16'b0000001110111110;
            15'd8829: log10_cal = 16'b0000001110111110;
            15'd8830: log10_cal = 16'b0000001110111110;
            15'd8831: log10_cal = 16'b0000001110111110;
            15'd8832: log10_cal = 16'b0000001110111110;
            15'd8833: log10_cal = 16'b0000001110111110;
            15'd8834: log10_cal = 16'b0000001110111110;
            15'd8835: log10_cal = 16'b0000001110111110;
            15'd8836: log10_cal = 16'b0000001110111110;
            15'd8837: log10_cal = 16'b0000001110111110;
            15'd8838: log10_cal = 16'b0000001110111110;
            15'd8839: log10_cal = 16'b0000001110111110;
            15'd8840: log10_cal = 16'b0000001110111110;
            15'd8841: log10_cal = 16'b0000001110111110;
            15'd8842: log10_cal = 16'b0000001110111110;
            15'd8843: log10_cal = 16'b0000001110111110;
            15'd8844: log10_cal = 16'b0000001110111110;
            15'd8845: log10_cal = 16'b0000001110111110;
            15'd8846: log10_cal = 16'b0000001110111110;
            15'd8847: log10_cal = 16'b0000001110111110;
            15'd8848: log10_cal = 16'b0000001110111111;
            15'd8849: log10_cal = 16'b0000001110111111;
            15'd8850: log10_cal = 16'b0000001110111111;
            15'd8851: log10_cal = 16'b0000001110111111;
            15'd8852: log10_cal = 16'b0000001110111111;
            15'd8853: log10_cal = 16'b0000001110111111;
            15'd8854: log10_cal = 16'b0000001110111111;
            15'd8855: log10_cal = 16'b0000001110111111;
            15'd8856: log10_cal = 16'b0000001110111111;
            15'd8857: log10_cal = 16'b0000001110111111;
            15'd8858: log10_cal = 16'b0000001110111111;
            15'd8859: log10_cal = 16'b0000001110111111;
            15'd8860: log10_cal = 16'b0000001110111111;
            15'd8861: log10_cal = 16'b0000001110111111;
            15'd8862: log10_cal = 16'b0000001110111111;
            15'd8863: log10_cal = 16'b0000001110111111;
            15'd8864: log10_cal = 16'b0000001110111111;
            15'd8865: log10_cal = 16'b0000001110111111;
            15'd8866: log10_cal = 16'b0000001110111111;
            15'd8867: log10_cal = 16'b0000001110111111;
            15'd8868: log10_cal = 16'b0000001111000000;
            15'd8869: log10_cal = 16'b0000001111000000;
            15'd8870: log10_cal = 16'b0000001111000000;
            15'd8871: log10_cal = 16'b0000001111000000;
            15'd8872: log10_cal = 16'b0000001111000000;
            15'd8873: log10_cal = 16'b0000001111000000;
            15'd8874: log10_cal = 16'b0000001111000000;
            15'd8875: log10_cal = 16'b0000001111000000;
            15'd8876: log10_cal = 16'b0000001111000000;
            15'd8877: log10_cal = 16'b0000001111000000;
            15'd8878: log10_cal = 16'b0000001111000000;
            15'd8879: log10_cal = 16'b0000001111000000;
            15'd8880: log10_cal = 16'b0000001111000000;
            15'd8881: log10_cal = 16'b0000001111000000;
            15'd8882: log10_cal = 16'b0000001111000000;
            15'd8883: log10_cal = 16'b0000001111000000;
            15'd8884: log10_cal = 16'b0000001111000000;
            15'd8885: log10_cal = 16'b0000001111000000;
            15'd8886: log10_cal = 16'b0000001111000000;
            15'd8887: log10_cal = 16'b0000001111000000;
            15'd8888: log10_cal = 16'b0000001111000001;
            15'd8889: log10_cal = 16'b0000001111000001;
            15'd8890: log10_cal = 16'b0000001111000001;
            15'd8891: log10_cal = 16'b0000001111000001;
            15'd8892: log10_cal = 16'b0000001111000001;
            15'd8893: log10_cal = 16'b0000001111000001;
            15'd8894: log10_cal = 16'b0000001111000001;
            15'd8895: log10_cal = 16'b0000001111000001;
            15'd8896: log10_cal = 16'b0000001111000001;
            15'd8897: log10_cal = 16'b0000001111000001;
            15'd8898: log10_cal = 16'b0000001111000001;
            15'd8899: log10_cal = 16'b0000001111000001;
            15'd8900: log10_cal = 16'b0000001111000001;
            15'd8901: log10_cal = 16'b0000001111000001;
            15'd8902: log10_cal = 16'b0000001111000001;
            15'd8903: log10_cal = 16'b0000001111000001;
            15'd8904: log10_cal = 16'b0000001111000001;
            15'd8905: log10_cal = 16'b0000001111000001;
            15'd8906: log10_cal = 16'b0000001111000001;
            15'd8907: log10_cal = 16'b0000001111000001;
            15'd8908: log10_cal = 16'b0000001111000010;
            15'd8909: log10_cal = 16'b0000001111000010;
            15'd8910: log10_cal = 16'b0000001111000010;
            15'd8911: log10_cal = 16'b0000001111000010;
            15'd8912: log10_cal = 16'b0000001111000010;
            15'd8913: log10_cal = 16'b0000001111000010;
            15'd8914: log10_cal = 16'b0000001111000010;
            15'd8915: log10_cal = 16'b0000001111000010;
            15'd8916: log10_cal = 16'b0000001111000010;
            15'd8917: log10_cal = 16'b0000001111000010;
            15'd8918: log10_cal = 16'b0000001111000010;
            15'd8919: log10_cal = 16'b0000001111000010;
            15'd8920: log10_cal = 16'b0000001111000010;
            15'd8921: log10_cal = 16'b0000001111000010;
            15'd8922: log10_cal = 16'b0000001111000010;
            15'd8923: log10_cal = 16'b0000001111000010;
            15'd8924: log10_cal = 16'b0000001111000010;
            15'd8925: log10_cal = 16'b0000001111000010;
            15'd8926: log10_cal = 16'b0000001111000010;
            15'd8927: log10_cal = 16'b0000001111000010;
            15'd8928: log10_cal = 16'b0000001111000011;
            15'd8929: log10_cal = 16'b0000001111000011;
            15'd8930: log10_cal = 16'b0000001111000011;
            15'd8931: log10_cal = 16'b0000001111000011;
            15'd8932: log10_cal = 16'b0000001111000011;
            15'd8933: log10_cal = 16'b0000001111000011;
            15'd8934: log10_cal = 16'b0000001111000011;
            15'd8935: log10_cal = 16'b0000001111000011;
            15'd8936: log10_cal = 16'b0000001111000011;
            15'd8937: log10_cal = 16'b0000001111000011;
            15'd8938: log10_cal = 16'b0000001111000011;
            15'd8939: log10_cal = 16'b0000001111000011;
            15'd8940: log10_cal = 16'b0000001111000011;
            15'd8941: log10_cal = 16'b0000001111000011;
            15'd8942: log10_cal = 16'b0000001111000011;
            15'd8943: log10_cal = 16'b0000001111000011;
            15'd8944: log10_cal = 16'b0000001111000011;
            15'd8945: log10_cal = 16'b0000001111000011;
            15'd8946: log10_cal = 16'b0000001111000011;
            15'd8947: log10_cal = 16'b0000001111000011;
            15'd8948: log10_cal = 16'b0000001111000100;
            15'd8949: log10_cal = 16'b0000001111000100;
            15'd8950: log10_cal = 16'b0000001111000100;
            15'd8951: log10_cal = 16'b0000001111000100;
            15'd8952: log10_cal = 16'b0000001111000100;
            15'd8953: log10_cal = 16'b0000001111000100;
            15'd8954: log10_cal = 16'b0000001111000100;
            15'd8955: log10_cal = 16'b0000001111000100;
            15'd8956: log10_cal = 16'b0000001111000100;
            15'd8957: log10_cal = 16'b0000001111000100;
            15'd8958: log10_cal = 16'b0000001111000100;
            15'd8959: log10_cal = 16'b0000001111000100;
            15'd8960: log10_cal = 16'b0000001111000100;
            15'd8961: log10_cal = 16'b0000001111000100;
            15'd8962: log10_cal = 16'b0000001111000100;
            15'd8963: log10_cal = 16'b0000001111000100;
            15'd8964: log10_cal = 16'b0000001111000100;
            15'd8965: log10_cal = 16'b0000001111000100;
            15'd8966: log10_cal = 16'b0000001111000100;
            15'd8967: log10_cal = 16'b0000001111000100;
            15'd8968: log10_cal = 16'b0000001111000101;
            15'd8969: log10_cal = 16'b0000001111000101;
            15'd8970: log10_cal = 16'b0000001111000101;
            15'd8971: log10_cal = 16'b0000001111000101;
            15'd8972: log10_cal = 16'b0000001111000101;
            15'd8973: log10_cal = 16'b0000001111000101;
            15'd8974: log10_cal = 16'b0000001111000101;
            15'd8975: log10_cal = 16'b0000001111000101;
            15'd8976: log10_cal = 16'b0000001111000101;
            15'd8977: log10_cal = 16'b0000001111000101;
            15'd8978: log10_cal = 16'b0000001111000101;
            15'd8979: log10_cal = 16'b0000001111000101;
            15'd8980: log10_cal = 16'b0000001111000101;
            15'd8981: log10_cal = 16'b0000001111000101;
            15'd8982: log10_cal = 16'b0000001111000101;
            15'd8983: log10_cal = 16'b0000001111000101;
            15'd8984: log10_cal = 16'b0000001111000101;
            15'd8985: log10_cal = 16'b0000001111000101;
            15'd8986: log10_cal = 16'b0000001111000101;
            15'd8987: log10_cal = 16'b0000001111000101;
            15'd8988: log10_cal = 16'b0000001111000110;
            15'd8989: log10_cal = 16'b0000001111000110;
            15'd8990: log10_cal = 16'b0000001111000110;
            15'd8991: log10_cal = 16'b0000001111000110;
            15'd8992: log10_cal = 16'b0000001111000110;
            15'd8993: log10_cal = 16'b0000001111000110;
            15'd8994: log10_cal = 16'b0000001111000110;
            15'd8995: log10_cal = 16'b0000001111000110;
            15'd8996: log10_cal = 16'b0000001111000110;
            15'd8997: log10_cal = 16'b0000001111000110;
            15'd8998: log10_cal = 16'b0000001111000110;
            15'd8999: log10_cal = 16'b0000001111000110;
            15'd9000: log10_cal = 16'b0000001111000110;
            15'd9001: log10_cal = 16'b0000001111000110;
            15'd9002: log10_cal = 16'b0000001111000110;
            15'd9003: log10_cal = 16'b0000001111000110;
            15'd9004: log10_cal = 16'b0000001111000110;
            15'd9005: log10_cal = 16'b0000001111000110;
            15'd9006: log10_cal = 16'b0000001111000110;
            15'd9007: log10_cal = 16'b0000001111000110;
            15'd9008: log10_cal = 16'b0000001111000110;
            15'd9009: log10_cal = 16'b0000001111000111;
            15'd9010: log10_cal = 16'b0000001111000111;
            15'd9011: log10_cal = 16'b0000001111000111;
            15'd9012: log10_cal = 16'b0000001111000111;
            15'd9013: log10_cal = 16'b0000001111000111;
            15'd9014: log10_cal = 16'b0000001111000111;
            15'd9015: log10_cal = 16'b0000001111000111;
            15'd9016: log10_cal = 16'b0000001111000111;
            15'd9017: log10_cal = 16'b0000001111000111;
            15'd9018: log10_cal = 16'b0000001111000111;
            15'd9019: log10_cal = 16'b0000001111000111;
            15'd9020: log10_cal = 16'b0000001111000111;
            15'd9021: log10_cal = 16'b0000001111000111;
            15'd9022: log10_cal = 16'b0000001111000111;
            15'd9023: log10_cal = 16'b0000001111000111;
            15'd9024: log10_cal = 16'b0000001111000111;
            15'd9025: log10_cal = 16'b0000001111000111;
            15'd9026: log10_cal = 16'b0000001111000111;
            15'd9027: log10_cal = 16'b0000001111000111;
            15'd9028: log10_cal = 16'b0000001111000111;
            15'd9029: log10_cal = 16'b0000001111001000;
            15'd9030: log10_cal = 16'b0000001111001000;
            15'd9031: log10_cal = 16'b0000001111001000;
            15'd9032: log10_cal = 16'b0000001111001000;
            15'd9033: log10_cal = 16'b0000001111001000;
            15'd9034: log10_cal = 16'b0000001111001000;
            15'd9035: log10_cal = 16'b0000001111001000;
            15'd9036: log10_cal = 16'b0000001111001000;
            15'd9037: log10_cal = 16'b0000001111001000;
            15'd9038: log10_cal = 16'b0000001111001000;
            15'd9039: log10_cal = 16'b0000001111001000;
            15'd9040: log10_cal = 16'b0000001111001000;
            15'd9041: log10_cal = 16'b0000001111001000;
            15'd9042: log10_cal = 16'b0000001111001000;
            15'd9043: log10_cal = 16'b0000001111001000;
            15'd9044: log10_cal = 16'b0000001111001000;
            15'd9045: log10_cal = 16'b0000001111001000;
            15'd9046: log10_cal = 16'b0000001111001000;
            15'd9047: log10_cal = 16'b0000001111001000;
            15'd9048: log10_cal = 16'b0000001111001000;
            15'd9049: log10_cal = 16'b0000001111001001;
            15'd9050: log10_cal = 16'b0000001111001001;
            15'd9051: log10_cal = 16'b0000001111001001;
            15'd9052: log10_cal = 16'b0000001111001001;
            15'd9053: log10_cal = 16'b0000001111001001;
            15'd9054: log10_cal = 16'b0000001111001001;
            15'd9055: log10_cal = 16'b0000001111001001;
            15'd9056: log10_cal = 16'b0000001111001001;
            15'd9057: log10_cal = 16'b0000001111001001;
            15'd9058: log10_cal = 16'b0000001111001001;
            15'd9059: log10_cal = 16'b0000001111001001;
            15'd9060: log10_cal = 16'b0000001111001001;
            15'd9061: log10_cal = 16'b0000001111001001;
            15'd9062: log10_cal = 16'b0000001111001001;
            15'd9063: log10_cal = 16'b0000001111001001;
            15'd9064: log10_cal = 16'b0000001111001001;
            15'd9065: log10_cal = 16'b0000001111001001;
            15'd9066: log10_cal = 16'b0000001111001001;
            15'd9067: log10_cal = 16'b0000001111001001;
            15'd9068: log10_cal = 16'b0000001111001001;
            15'd9069: log10_cal = 16'b0000001111001001;
            15'd9070: log10_cal = 16'b0000001111001010;
            15'd9071: log10_cal = 16'b0000001111001010;
            15'd9072: log10_cal = 16'b0000001111001010;
            15'd9073: log10_cal = 16'b0000001111001010;
            15'd9074: log10_cal = 16'b0000001111001010;
            15'd9075: log10_cal = 16'b0000001111001010;
            15'd9076: log10_cal = 16'b0000001111001010;
            15'd9077: log10_cal = 16'b0000001111001010;
            15'd9078: log10_cal = 16'b0000001111001010;
            15'd9079: log10_cal = 16'b0000001111001010;
            15'd9080: log10_cal = 16'b0000001111001010;
            15'd9081: log10_cal = 16'b0000001111001010;
            15'd9082: log10_cal = 16'b0000001111001010;
            15'd9083: log10_cal = 16'b0000001111001010;
            15'd9084: log10_cal = 16'b0000001111001010;
            15'd9085: log10_cal = 16'b0000001111001010;
            15'd9086: log10_cal = 16'b0000001111001010;
            15'd9087: log10_cal = 16'b0000001111001010;
            15'd9088: log10_cal = 16'b0000001111001010;
            15'd9089: log10_cal = 16'b0000001111001010;
            15'd9090: log10_cal = 16'b0000001111001011;
            15'd9091: log10_cal = 16'b0000001111001011;
            15'd9092: log10_cal = 16'b0000001111001011;
            15'd9093: log10_cal = 16'b0000001111001011;
            15'd9094: log10_cal = 16'b0000001111001011;
            15'd9095: log10_cal = 16'b0000001111001011;
            15'd9096: log10_cal = 16'b0000001111001011;
            15'd9097: log10_cal = 16'b0000001111001011;
            15'd9098: log10_cal = 16'b0000001111001011;
            15'd9099: log10_cal = 16'b0000001111001011;
            15'd9100: log10_cal = 16'b0000001111001011;
            15'd9101: log10_cal = 16'b0000001111001011;
            15'd9102: log10_cal = 16'b0000001111001011;
            15'd9103: log10_cal = 16'b0000001111001011;
            15'd9104: log10_cal = 16'b0000001111001011;
            15'd9105: log10_cal = 16'b0000001111001011;
            15'd9106: log10_cal = 16'b0000001111001011;
            15'd9107: log10_cal = 16'b0000001111001011;
            15'd9108: log10_cal = 16'b0000001111001011;
            15'd9109: log10_cal = 16'b0000001111001011;
            15'd9110: log10_cal = 16'b0000001111001011;
            15'd9111: log10_cal = 16'b0000001111001100;
            15'd9112: log10_cal = 16'b0000001111001100;
            15'd9113: log10_cal = 16'b0000001111001100;
            15'd9114: log10_cal = 16'b0000001111001100;
            15'd9115: log10_cal = 16'b0000001111001100;
            15'd9116: log10_cal = 16'b0000001111001100;
            15'd9117: log10_cal = 16'b0000001111001100;
            15'd9118: log10_cal = 16'b0000001111001100;
            15'd9119: log10_cal = 16'b0000001111001100;
            15'd9120: log10_cal = 16'b0000001111001100;
            15'd9121: log10_cal = 16'b0000001111001100;
            15'd9122: log10_cal = 16'b0000001111001100;
            15'd9123: log10_cal = 16'b0000001111001100;
            15'd9124: log10_cal = 16'b0000001111001100;
            15'd9125: log10_cal = 16'b0000001111001100;
            15'd9126: log10_cal = 16'b0000001111001100;
            15'd9127: log10_cal = 16'b0000001111001100;
            15'd9128: log10_cal = 16'b0000001111001100;
            15'd9129: log10_cal = 16'b0000001111001100;
            15'd9130: log10_cal = 16'b0000001111001100;
            15'd9131: log10_cal = 16'b0000001111001101;
            15'd9132: log10_cal = 16'b0000001111001101;
            15'd9133: log10_cal = 16'b0000001111001101;
            15'd9134: log10_cal = 16'b0000001111001101;
            15'd9135: log10_cal = 16'b0000001111001101;
            15'd9136: log10_cal = 16'b0000001111001101;
            15'd9137: log10_cal = 16'b0000001111001101;
            15'd9138: log10_cal = 16'b0000001111001101;
            15'd9139: log10_cal = 16'b0000001111001101;
            15'd9140: log10_cal = 16'b0000001111001101;
            15'd9141: log10_cal = 16'b0000001111001101;
            15'd9142: log10_cal = 16'b0000001111001101;
            15'd9143: log10_cal = 16'b0000001111001101;
            15'd9144: log10_cal = 16'b0000001111001101;
            15'd9145: log10_cal = 16'b0000001111001101;
            15'd9146: log10_cal = 16'b0000001111001101;
            15'd9147: log10_cal = 16'b0000001111001101;
            15'd9148: log10_cal = 16'b0000001111001101;
            15'd9149: log10_cal = 16'b0000001111001101;
            15'd9150: log10_cal = 16'b0000001111001101;
            15'd9151: log10_cal = 16'b0000001111001101;
            15'd9152: log10_cal = 16'b0000001111001110;
            15'd9153: log10_cal = 16'b0000001111001110;
            15'd9154: log10_cal = 16'b0000001111001110;
            15'd9155: log10_cal = 16'b0000001111001110;
            15'd9156: log10_cal = 16'b0000001111001110;
            15'd9157: log10_cal = 16'b0000001111001110;
            15'd9158: log10_cal = 16'b0000001111001110;
            15'd9159: log10_cal = 16'b0000001111001110;
            15'd9160: log10_cal = 16'b0000001111001110;
            15'd9161: log10_cal = 16'b0000001111001110;
            15'd9162: log10_cal = 16'b0000001111001110;
            15'd9163: log10_cal = 16'b0000001111001110;
            15'd9164: log10_cal = 16'b0000001111001110;
            15'd9165: log10_cal = 16'b0000001111001110;
            15'd9166: log10_cal = 16'b0000001111001110;
            15'd9167: log10_cal = 16'b0000001111001110;
            15'd9168: log10_cal = 16'b0000001111001110;
            15'd9169: log10_cal = 16'b0000001111001110;
            15'd9170: log10_cal = 16'b0000001111001110;
            15'd9171: log10_cal = 16'b0000001111001110;
            15'd9172: log10_cal = 16'b0000001111001111;
            15'd9173: log10_cal = 16'b0000001111001111;
            15'd9174: log10_cal = 16'b0000001111001111;
            15'd9175: log10_cal = 16'b0000001111001111;
            15'd9176: log10_cal = 16'b0000001111001111;
            15'd9177: log10_cal = 16'b0000001111001111;
            15'd9178: log10_cal = 16'b0000001111001111;
            15'd9179: log10_cal = 16'b0000001111001111;
            15'd9180: log10_cal = 16'b0000001111001111;
            15'd9181: log10_cal = 16'b0000001111001111;
            15'd9182: log10_cal = 16'b0000001111001111;
            15'd9183: log10_cal = 16'b0000001111001111;
            15'd9184: log10_cal = 16'b0000001111001111;
            15'd9185: log10_cal = 16'b0000001111001111;
            15'd9186: log10_cal = 16'b0000001111001111;
            15'd9187: log10_cal = 16'b0000001111001111;
            15'd9188: log10_cal = 16'b0000001111001111;
            15'd9189: log10_cal = 16'b0000001111001111;
            15'd9190: log10_cal = 16'b0000001111001111;
            15'd9191: log10_cal = 16'b0000001111001111;
            15'd9192: log10_cal = 16'b0000001111001111;
            15'd9193: log10_cal = 16'b0000001111010000;
            15'd9194: log10_cal = 16'b0000001111010000;
            15'd9195: log10_cal = 16'b0000001111010000;
            15'd9196: log10_cal = 16'b0000001111010000;
            15'd9197: log10_cal = 16'b0000001111010000;
            15'd9198: log10_cal = 16'b0000001111010000;
            15'd9199: log10_cal = 16'b0000001111010000;
            15'd9200: log10_cal = 16'b0000001111010000;
            15'd9201: log10_cal = 16'b0000001111010000;
            15'd9202: log10_cal = 16'b0000001111010000;
            15'd9203: log10_cal = 16'b0000001111010000;
            15'd9204: log10_cal = 16'b0000001111010000;
            15'd9205: log10_cal = 16'b0000001111010000;
            15'd9206: log10_cal = 16'b0000001111010000;
            15'd9207: log10_cal = 16'b0000001111010000;
            15'd9208: log10_cal = 16'b0000001111010000;
            15'd9209: log10_cal = 16'b0000001111010000;
            15'd9210: log10_cal = 16'b0000001111010000;
            15'd9211: log10_cal = 16'b0000001111010000;
            15'd9212: log10_cal = 16'b0000001111010000;
            15'd9213: log10_cal = 16'b0000001111010000;
            15'd9214: log10_cal = 16'b0000001111010001;
            15'd9215: log10_cal = 16'b0000001111010001;
            15'd9216: log10_cal = 16'b0000001111010001;
            15'd9217: log10_cal = 16'b0000001111010001;
            15'd9218: log10_cal = 16'b0000001111010001;
            15'd9219: log10_cal = 16'b0000001111010001;
            15'd9220: log10_cal = 16'b0000001111010001;
            15'd9221: log10_cal = 16'b0000001111010001;
            15'd9222: log10_cal = 16'b0000001111010001;
            15'd9223: log10_cal = 16'b0000001111010001;
            15'd9224: log10_cal = 16'b0000001111010001;
            15'd9225: log10_cal = 16'b0000001111010001;
            15'd9226: log10_cal = 16'b0000001111010001;
            15'd9227: log10_cal = 16'b0000001111010001;
            15'd9228: log10_cal = 16'b0000001111010001;
            15'd9229: log10_cal = 16'b0000001111010001;
            15'd9230: log10_cal = 16'b0000001111010001;
            15'd9231: log10_cal = 16'b0000001111010001;
            15'd9232: log10_cal = 16'b0000001111010001;
            15'd9233: log10_cal = 16'b0000001111010001;
            15'd9234: log10_cal = 16'b0000001111010010;
            15'd9235: log10_cal = 16'b0000001111010010;
            15'd9236: log10_cal = 16'b0000001111010010;
            15'd9237: log10_cal = 16'b0000001111010010;
            15'd9238: log10_cal = 16'b0000001111010010;
            15'd9239: log10_cal = 16'b0000001111010010;
            15'd9240: log10_cal = 16'b0000001111010010;
            15'd9241: log10_cal = 16'b0000001111010010;
            15'd9242: log10_cal = 16'b0000001111010010;
            15'd9243: log10_cal = 16'b0000001111010010;
            15'd9244: log10_cal = 16'b0000001111010010;
            15'd9245: log10_cal = 16'b0000001111010010;
            15'd9246: log10_cal = 16'b0000001111010010;
            15'd9247: log10_cal = 16'b0000001111010010;
            15'd9248: log10_cal = 16'b0000001111010010;
            15'd9249: log10_cal = 16'b0000001111010010;
            15'd9250: log10_cal = 16'b0000001111010010;
            15'd9251: log10_cal = 16'b0000001111010010;
            15'd9252: log10_cal = 16'b0000001111010010;
            15'd9253: log10_cal = 16'b0000001111010010;
            15'd9254: log10_cal = 16'b0000001111010010;
            15'd9255: log10_cal = 16'b0000001111010011;
            15'd9256: log10_cal = 16'b0000001111010011;
            15'd9257: log10_cal = 16'b0000001111010011;
            15'd9258: log10_cal = 16'b0000001111010011;
            15'd9259: log10_cal = 16'b0000001111010011;
            15'd9260: log10_cal = 16'b0000001111010011;
            15'd9261: log10_cal = 16'b0000001111010011;
            15'd9262: log10_cal = 16'b0000001111010011;
            15'd9263: log10_cal = 16'b0000001111010011;
            15'd9264: log10_cal = 16'b0000001111010011;
            15'd9265: log10_cal = 16'b0000001111010011;
            15'd9266: log10_cal = 16'b0000001111010011;
            15'd9267: log10_cal = 16'b0000001111010011;
            15'd9268: log10_cal = 16'b0000001111010011;
            15'd9269: log10_cal = 16'b0000001111010011;
            15'd9270: log10_cal = 16'b0000001111010011;
            15'd9271: log10_cal = 16'b0000001111010011;
            15'd9272: log10_cal = 16'b0000001111010011;
            15'd9273: log10_cal = 16'b0000001111010011;
            15'd9274: log10_cal = 16'b0000001111010011;
            15'd9275: log10_cal = 16'b0000001111010011;
            15'd9276: log10_cal = 16'b0000001111010100;
            15'd9277: log10_cal = 16'b0000001111010100;
            15'd9278: log10_cal = 16'b0000001111010100;
            15'd9279: log10_cal = 16'b0000001111010100;
            15'd9280: log10_cal = 16'b0000001111010100;
            15'd9281: log10_cal = 16'b0000001111010100;
            15'd9282: log10_cal = 16'b0000001111010100;
            15'd9283: log10_cal = 16'b0000001111010100;
            15'd9284: log10_cal = 16'b0000001111010100;
            15'd9285: log10_cal = 16'b0000001111010100;
            15'd9286: log10_cal = 16'b0000001111010100;
            15'd9287: log10_cal = 16'b0000001111010100;
            15'd9288: log10_cal = 16'b0000001111010100;
            15'd9289: log10_cal = 16'b0000001111010100;
            15'd9290: log10_cal = 16'b0000001111010100;
            15'd9291: log10_cal = 16'b0000001111010100;
            15'd9292: log10_cal = 16'b0000001111010100;
            15'd9293: log10_cal = 16'b0000001111010100;
            15'd9294: log10_cal = 16'b0000001111010100;
            15'd9295: log10_cal = 16'b0000001111010100;
            15'd9296: log10_cal = 16'b0000001111010100;
            15'd9297: log10_cal = 16'b0000001111010101;
            15'd9298: log10_cal = 16'b0000001111010101;
            15'd9299: log10_cal = 16'b0000001111010101;
            15'd9300: log10_cal = 16'b0000001111010101;
            15'd9301: log10_cal = 16'b0000001111010101;
            15'd9302: log10_cal = 16'b0000001111010101;
            15'd9303: log10_cal = 16'b0000001111010101;
            15'd9304: log10_cal = 16'b0000001111010101;
            15'd9305: log10_cal = 16'b0000001111010101;
            15'd9306: log10_cal = 16'b0000001111010101;
            15'd9307: log10_cal = 16'b0000001111010101;
            15'd9308: log10_cal = 16'b0000001111010101;
            15'd9309: log10_cal = 16'b0000001111010101;
            15'd9310: log10_cal = 16'b0000001111010101;
            15'd9311: log10_cal = 16'b0000001111010101;
            15'd9312: log10_cal = 16'b0000001111010101;
            15'd9313: log10_cal = 16'b0000001111010101;
            15'd9314: log10_cal = 16'b0000001111010101;
            15'd9315: log10_cal = 16'b0000001111010101;
            15'd9316: log10_cal = 16'b0000001111010101;
            15'd9317: log10_cal = 16'b0000001111010101;
            15'd9318: log10_cal = 16'b0000001111010110;
            15'd9319: log10_cal = 16'b0000001111010110;
            15'd9320: log10_cal = 16'b0000001111010110;
            15'd9321: log10_cal = 16'b0000001111010110;
            15'd9322: log10_cal = 16'b0000001111010110;
            15'd9323: log10_cal = 16'b0000001111010110;
            15'd9324: log10_cal = 16'b0000001111010110;
            15'd9325: log10_cal = 16'b0000001111010110;
            15'd9326: log10_cal = 16'b0000001111010110;
            15'd9327: log10_cal = 16'b0000001111010110;
            15'd9328: log10_cal = 16'b0000001111010110;
            15'd9329: log10_cal = 16'b0000001111010110;
            15'd9330: log10_cal = 16'b0000001111010110;
            15'd9331: log10_cal = 16'b0000001111010110;
            15'd9332: log10_cal = 16'b0000001111010110;
            15'd9333: log10_cal = 16'b0000001111010110;
            15'd9334: log10_cal = 16'b0000001111010110;
            15'd9335: log10_cal = 16'b0000001111010110;
            15'd9336: log10_cal = 16'b0000001111010110;
            15'd9337: log10_cal = 16'b0000001111010110;
            15'd9338: log10_cal = 16'b0000001111010110;
            15'd9339: log10_cal = 16'b0000001111010111;
            15'd9340: log10_cal = 16'b0000001111010111;
            15'd9341: log10_cal = 16'b0000001111010111;
            15'd9342: log10_cal = 16'b0000001111010111;
            15'd9343: log10_cal = 16'b0000001111010111;
            15'd9344: log10_cal = 16'b0000001111010111;
            15'd9345: log10_cal = 16'b0000001111010111;
            15'd9346: log10_cal = 16'b0000001111010111;
            15'd9347: log10_cal = 16'b0000001111010111;
            15'd9348: log10_cal = 16'b0000001111010111;
            15'd9349: log10_cal = 16'b0000001111010111;
            15'd9350: log10_cal = 16'b0000001111010111;
            15'd9351: log10_cal = 16'b0000001111010111;
            15'd9352: log10_cal = 16'b0000001111010111;
            15'd9353: log10_cal = 16'b0000001111010111;
            15'd9354: log10_cal = 16'b0000001111010111;
            15'd9355: log10_cal = 16'b0000001111010111;
            15'd9356: log10_cal = 16'b0000001111010111;
            15'd9357: log10_cal = 16'b0000001111010111;
            15'd9358: log10_cal = 16'b0000001111010111;
            15'd9359: log10_cal = 16'b0000001111010111;
            15'd9360: log10_cal = 16'b0000001111011000;
            15'd9361: log10_cal = 16'b0000001111011000;
            15'd9362: log10_cal = 16'b0000001111011000;
            15'd9363: log10_cal = 16'b0000001111011000;
            15'd9364: log10_cal = 16'b0000001111011000;
            15'd9365: log10_cal = 16'b0000001111011000;
            15'd9366: log10_cal = 16'b0000001111011000;
            15'd9367: log10_cal = 16'b0000001111011000;
            15'd9368: log10_cal = 16'b0000001111011000;
            15'd9369: log10_cal = 16'b0000001111011000;
            15'd9370: log10_cal = 16'b0000001111011000;
            15'd9371: log10_cal = 16'b0000001111011000;
            15'd9372: log10_cal = 16'b0000001111011000;
            15'd9373: log10_cal = 16'b0000001111011000;
            15'd9374: log10_cal = 16'b0000001111011000;
            15'd9375: log10_cal = 16'b0000001111011000;
            15'd9376: log10_cal = 16'b0000001111011000;
            15'd9377: log10_cal = 16'b0000001111011000;
            15'd9378: log10_cal = 16'b0000001111011000;
            15'd9379: log10_cal = 16'b0000001111011000;
            15'd9380: log10_cal = 16'b0000001111011000;
            15'd9381: log10_cal = 16'b0000001111011001;
            15'd9382: log10_cal = 16'b0000001111011001;
            15'd9383: log10_cal = 16'b0000001111011001;
            15'd9384: log10_cal = 16'b0000001111011001;
            15'd9385: log10_cal = 16'b0000001111011001;
            15'd9386: log10_cal = 16'b0000001111011001;
            15'd9387: log10_cal = 16'b0000001111011001;
            15'd9388: log10_cal = 16'b0000001111011001;
            15'd9389: log10_cal = 16'b0000001111011001;
            15'd9390: log10_cal = 16'b0000001111011001;
            15'd9391: log10_cal = 16'b0000001111011001;
            15'd9392: log10_cal = 16'b0000001111011001;
            15'd9393: log10_cal = 16'b0000001111011001;
            15'd9394: log10_cal = 16'b0000001111011001;
            15'd9395: log10_cal = 16'b0000001111011001;
            15'd9396: log10_cal = 16'b0000001111011001;
            15'd9397: log10_cal = 16'b0000001111011001;
            15'd9398: log10_cal = 16'b0000001111011001;
            15'd9399: log10_cal = 16'b0000001111011001;
            15'd9400: log10_cal = 16'b0000001111011001;
            15'd9401: log10_cal = 16'b0000001111011001;
            15'd9402: log10_cal = 16'b0000001111011010;
            15'd9403: log10_cal = 16'b0000001111011010;
            15'd9404: log10_cal = 16'b0000001111011010;
            15'd9405: log10_cal = 16'b0000001111011010;
            15'd9406: log10_cal = 16'b0000001111011010;
            15'd9407: log10_cal = 16'b0000001111011010;
            15'd9408: log10_cal = 16'b0000001111011010;
            15'd9409: log10_cal = 16'b0000001111011010;
            15'd9410: log10_cal = 16'b0000001111011010;
            15'd9411: log10_cal = 16'b0000001111011010;
            15'd9412: log10_cal = 16'b0000001111011010;
            15'd9413: log10_cal = 16'b0000001111011010;
            15'd9414: log10_cal = 16'b0000001111011010;
            15'd9415: log10_cal = 16'b0000001111011010;
            15'd9416: log10_cal = 16'b0000001111011010;
            15'd9417: log10_cal = 16'b0000001111011010;
            15'd9418: log10_cal = 16'b0000001111011010;
            15'd9419: log10_cal = 16'b0000001111011010;
            15'd9420: log10_cal = 16'b0000001111011010;
            15'd9421: log10_cal = 16'b0000001111011010;
            15'd9422: log10_cal = 16'b0000001111011010;
            15'd9423: log10_cal = 16'b0000001111011011;
            15'd9424: log10_cal = 16'b0000001111011011;
            15'd9425: log10_cal = 16'b0000001111011011;
            15'd9426: log10_cal = 16'b0000001111011011;
            15'd9427: log10_cal = 16'b0000001111011011;
            15'd9428: log10_cal = 16'b0000001111011011;
            15'd9429: log10_cal = 16'b0000001111011011;
            15'd9430: log10_cal = 16'b0000001111011011;
            15'd9431: log10_cal = 16'b0000001111011011;
            15'd9432: log10_cal = 16'b0000001111011011;
            15'd9433: log10_cal = 16'b0000001111011011;
            15'd9434: log10_cal = 16'b0000001111011011;
            15'd9435: log10_cal = 16'b0000001111011011;
            15'd9436: log10_cal = 16'b0000001111011011;
            15'd9437: log10_cal = 16'b0000001111011011;
            15'd9438: log10_cal = 16'b0000001111011011;
            15'd9439: log10_cal = 16'b0000001111011011;
            15'd9440: log10_cal = 16'b0000001111011011;
            15'd9441: log10_cal = 16'b0000001111011011;
            15'd9442: log10_cal = 16'b0000001111011011;
            15'd9443: log10_cal = 16'b0000001111011011;
            15'd9444: log10_cal = 16'b0000001111011100;
            15'd9445: log10_cal = 16'b0000001111011100;
            15'd9446: log10_cal = 16'b0000001111011100;
            15'd9447: log10_cal = 16'b0000001111011100;
            15'd9448: log10_cal = 16'b0000001111011100;
            15'd9449: log10_cal = 16'b0000001111011100;
            15'd9450: log10_cal = 16'b0000001111011100;
            15'd9451: log10_cal = 16'b0000001111011100;
            15'd9452: log10_cal = 16'b0000001111011100;
            15'd9453: log10_cal = 16'b0000001111011100;
            15'd9454: log10_cal = 16'b0000001111011100;
            15'd9455: log10_cal = 16'b0000001111011100;
            15'd9456: log10_cal = 16'b0000001111011100;
            15'd9457: log10_cal = 16'b0000001111011100;
            15'd9458: log10_cal = 16'b0000001111011100;
            15'd9459: log10_cal = 16'b0000001111011100;
            15'd9460: log10_cal = 16'b0000001111011100;
            15'd9461: log10_cal = 16'b0000001111011100;
            15'd9462: log10_cal = 16'b0000001111011100;
            15'd9463: log10_cal = 16'b0000001111011100;
            15'd9464: log10_cal = 16'b0000001111011100;
            15'd9465: log10_cal = 16'b0000001111011101;
            15'd9466: log10_cal = 16'b0000001111011101;
            15'd9467: log10_cal = 16'b0000001111011101;
            15'd9468: log10_cal = 16'b0000001111011101;
            15'd9469: log10_cal = 16'b0000001111011101;
            15'd9470: log10_cal = 16'b0000001111011101;
            15'd9471: log10_cal = 16'b0000001111011101;
            15'd9472: log10_cal = 16'b0000001111011101;
            15'd9473: log10_cal = 16'b0000001111011101;
            15'd9474: log10_cal = 16'b0000001111011101;
            15'd9475: log10_cal = 16'b0000001111011101;
            15'd9476: log10_cal = 16'b0000001111011101;
            15'd9477: log10_cal = 16'b0000001111011101;
            15'd9478: log10_cal = 16'b0000001111011101;
            15'd9479: log10_cal = 16'b0000001111011101;
            15'd9480: log10_cal = 16'b0000001111011101;
            15'd9481: log10_cal = 16'b0000001111011101;
            15'd9482: log10_cal = 16'b0000001111011101;
            15'd9483: log10_cal = 16'b0000001111011101;
            15'd9484: log10_cal = 16'b0000001111011101;
            15'd9485: log10_cal = 16'b0000001111011101;
            15'd9486: log10_cal = 16'b0000001111011101;
            15'd9487: log10_cal = 16'b0000001111011110;
            15'd9488: log10_cal = 16'b0000001111011110;
            15'd9489: log10_cal = 16'b0000001111011110;
            15'd9490: log10_cal = 16'b0000001111011110;
            15'd9491: log10_cal = 16'b0000001111011110;
            15'd9492: log10_cal = 16'b0000001111011110;
            15'd9493: log10_cal = 16'b0000001111011110;
            15'd9494: log10_cal = 16'b0000001111011110;
            15'd9495: log10_cal = 16'b0000001111011110;
            15'd9496: log10_cal = 16'b0000001111011110;
            15'd9497: log10_cal = 16'b0000001111011110;
            15'd9498: log10_cal = 16'b0000001111011110;
            15'd9499: log10_cal = 16'b0000001111011110;
            15'd9500: log10_cal = 16'b0000001111011110;
            15'd9501: log10_cal = 16'b0000001111011110;
            15'd9502: log10_cal = 16'b0000001111011110;
            15'd9503: log10_cal = 16'b0000001111011110;
            15'd9504: log10_cal = 16'b0000001111011110;
            15'd9505: log10_cal = 16'b0000001111011110;
            15'd9506: log10_cal = 16'b0000001111011110;
            15'd9507: log10_cal = 16'b0000001111011110;
            15'd9508: log10_cal = 16'b0000001111011111;
            15'd9509: log10_cal = 16'b0000001111011111;
            15'd9510: log10_cal = 16'b0000001111011111;
            15'd9511: log10_cal = 16'b0000001111011111;
            15'd9512: log10_cal = 16'b0000001111011111;
            15'd9513: log10_cal = 16'b0000001111011111;
            15'd9514: log10_cal = 16'b0000001111011111;
            15'd9515: log10_cal = 16'b0000001111011111;
            15'd9516: log10_cal = 16'b0000001111011111;
            15'd9517: log10_cal = 16'b0000001111011111;
            15'd9518: log10_cal = 16'b0000001111011111;
            15'd9519: log10_cal = 16'b0000001111011111;
            15'd9520: log10_cal = 16'b0000001111011111;
            15'd9521: log10_cal = 16'b0000001111011111;
            15'd9522: log10_cal = 16'b0000001111011111;
            15'd9523: log10_cal = 16'b0000001111011111;
            15'd9524: log10_cal = 16'b0000001111011111;
            15'd9525: log10_cal = 16'b0000001111011111;
            15'd9526: log10_cal = 16'b0000001111011111;
            15'd9527: log10_cal = 16'b0000001111011111;
            15'd9528: log10_cal = 16'b0000001111011111;
            15'd9529: log10_cal = 16'b0000001111011111;
            15'd9530: log10_cal = 16'b0000001111100000;
            15'd9531: log10_cal = 16'b0000001111100000;
            15'd9532: log10_cal = 16'b0000001111100000;
            15'd9533: log10_cal = 16'b0000001111100000;
            15'd9534: log10_cal = 16'b0000001111100000;
            15'd9535: log10_cal = 16'b0000001111100000;
            15'd9536: log10_cal = 16'b0000001111100000;
            15'd9537: log10_cal = 16'b0000001111100000;
            15'd9538: log10_cal = 16'b0000001111100000;
            15'd9539: log10_cal = 16'b0000001111100000;
            15'd9540: log10_cal = 16'b0000001111100000;
            15'd9541: log10_cal = 16'b0000001111100000;
            15'd9542: log10_cal = 16'b0000001111100000;
            15'd9543: log10_cal = 16'b0000001111100000;
            15'd9544: log10_cal = 16'b0000001111100000;
            15'd9545: log10_cal = 16'b0000001111100000;
            15'd9546: log10_cal = 16'b0000001111100000;
            15'd9547: log10_cal = 16'b0000001111100000;
            15'd9548: log10_cal = 16'b0000001111100000;
            15'd9549: log10_cal = 16'b0000001111100000;
            15'd9550: log10_cal = 16'b0000001111100000;
            15'd9551: log10_cal = 16'b0000001111100001;
            15'd9552: log10_cal = 16'b0000001111100001;
            15'd9553: log10_cal = 16'b0000001111100001;
            15'd9554: log10_cal = 16'b0000001111100001;
            15'd9555: log10_cal = 16'b0000001111100001;
            15'd9556: log10_cal = 16'b0000001111100001;
            15'd9557: log10_cal = 16'b0000001111100001;
            15'd9558: log10_cal = 16'b0000001111100001;
            15'd9559: log10_cal = 16'b0000001111100001;
            15'd9560: log10_cal = 16'b0000001111100001;
            15'd9561: log10_cal = 16'b0000001111100001;
            15'd9562: log10_cal = 16'b0000001111100001;
            15'd9563: log10_cal = 16'b0000001111100001;
            15'd9564: log10_cal = 16'b0000001111100001;
            15'd9565: log10_cal = 16'b0000001111100001;
            15'd9566: log10_cal = 16'b0000001111100001;
            15'd9567: log10_cal = 16'b0000001111100001;
            15'd9568: log10_cal = 16'b0000001111100001;
            15'd9569: log10_cal = 16'b0000001111100001;
            15'd9570: log10_cal = 16'b0000001111100001;
            15'd9571: log10_cal = 16'b0000001111100001;
            15'd9572: log10_cal = 16'b0000001111100001;
            15'd9573: log10_cal = 16'b0000001111100010;
            15'd9574: log10_cal = 16'b0000001111100010;
            15'd9575: log10_cal = 16'b0000001111100010;
            15'd9576: log10_cal = 16'b0000001111100010;
            15'd9577: log10_cal = 16'b0000001111100010;
            15'd9578: log10_cal = 16'b0000001111100010;
            15'd9579: log10_cal = 16'b0000001111100010;
            15'd9580: log10_cal = 16'b0000001111100010;
            15'd9581: log10_cal = 16'b0000001111100010;
            15'd9582: log10_cal = 16'b0000001111100010;
            15'd9583: log10_cal = 16'b0000001111100010;
            15'd9584: log10_cal = 16'b0000001111100010;
            15'd9585: log10_cal = 16'b0000001111100010;
            15'd9586: log10_cal = 16'b0000001111100010;
            15'd9587: log10_cal = 16'b0000001111100010;
            15'd9588: log10_cal = 16'b0000001111100010;
            15'd9589: log10_cal = 16'b0000001111100010;
            15'd9590: log10_cal = 16'b0000001111100010;
            15'd9591: log10_cal = 16'b0000001111100010;
            15'd9592: log10_cal = 16'b0000001111100010;
            15'd9593: log10_cal = 16'b0000001111100010;
            15'd9594: log10_cal = 16'b0000001111100011;
            15'd9595: log10_cal = 16'b0000001111100011;
            15'd9596: log10_cal = 16'b0000001111100011;
            15'd9597: log10_cal = 16'b0000001111100011;
            15'd9598: log10_cal = 16'b0000001111100011;
            15'd9599: log10_cal = 16'b0000001111100011;
            15'd9600: log10_cal = 16'b0000001111100011;
            15'd9601: log10_cal = 16'b0000001111100011;
            15'd9602: log10_cal = 16'b0000001111100011;
            15'd9603: log10_cal = 16'b0000001111100011;
            15'd9604: log10_cal = 16'b0000001111100011;
            15'd9605: log10_cal = 16'b0000001111100011;
            15'd9606: log10_cal = 16'b0000001111100011;
            15'd9607: log10_cal = 16'b0000001111100011;
            15'd9608: log10_cal = 16'b0000001111100011;
            15'd9609: log10_cal = 16'b0000001111100011;
            15'd9610: log10_cal = 16'b0000001111100011;
            15'd9611: log10_cal = 16'b0000001111100011;
            15'd9612: log10_cal = 16'b0000001111100011;
            15'd9613: log10_cal = 16'b0000001111100011;
            15'd9614: log10_cal = 16'b0000001111100011;
            15'd9615: log10_cal = 16'b0000001111100011;
            15'd9616: log10_cal = 16'b0000001111100100;
            15'd9617: log10_cal = 16'b0000001111100100;
            15'd9618: log10_cal = 16'b0000001111100100;
            15'd9619: log10_cal = 16'b0000001111100100;
            15'd9620: log10_cal = 16'b0000001111100100;
            15'd9621: log10_cal = 16'b0000001111100100;
            15'd9622: log10_cal = 16'b0000001111100100;
            15'd9623: log10_cal = 16'b0000001111100100;
            15'd9624: log10_cal = 16'b0000001111100100;
            15'd9625: log10_cal = 16'b0000001111100100;
            15'd9626: log10_cal = 16'b0000001111100100;
            15'd9627: log10_cal = 16'b0000001111100100;
            15'd9628: log10_cal = 16'b0000001111100100;
            15'd9629: log10_cal = 16'b0000001111100100;
            15'd9630: log10_cal = 16'b0000001111100100;
            15'd9631: log10_cal = 16'b0000001111100100;
            15'd9632: log10_cal = 16'b0000001111100100;
            15'd9633: log10_cal = 16'b0000001111100100;
            15'd9634: log10_cal = 16'b0000001111100100;
            15'd9635: log10_cal = 16'b0000001111100100;
            15'd9636: log10_cal = 16'b0000001111100100;
            15'd9637: log10_cal = 16'b0000001111100101;
            15'd9638: log10_cal = 16'b0000001111100101;
            15'd9639: log10_cal = 16'b0000001111100101;
            15'd9640: log10_cal = 16'b0000001111100101;
            15'd9641: log10_cal = 16'b0000001111100101;
            15'd9642: log10_cal = 16'b0000001111100101;
            15'd9643: log10_cal = 16'b0000001111100101;
            15'd9644: log10_cal = 16'b0000001111100101;
            15'd9645: log10_cal = 16'b0000001111100101;
            15'd9646: log10_cal = 16'b0000001111100101;
            15'd9647: log10_cal = 16'b0000001111100101;
            15'd9648: log10_cal = 16'b0000001111100101;
            15'd9649: log10_cal = 16'b0000001111100101;
            15'd9650: log10_cal = 16'b0000001111100101;
            15'd9651: log10_cal = 16'b0000001111100101;
            15'd9652: log10_cal = 16'b0000001111100101;
            15'd9653: log10_cal = 16'b0000001111100101;
            15'd9654: log10_cal = 16'b0000001111100101;
            15'd9655: log10_cal = 16'b0000001111100101;
            15'd9656: log10_cal = 16'b0000001111100101;
            15'd9657: log10_cal = 16'b0000001111100101;
            15'd9658: log10_cal = 16'b0000001111100101;
            15'd9659: log10_cal = 16'b0000001111100110;
            15'd9660: log10_cal = 16'b0000001111100110;
            15'd9661: log10_cal = 16'b0000001111100110;
            15'd9662: log10_cal = 16'b0000001111100110;
            15'd9663: log10_cal = 16'b0000001111100110;
            15'd9664: log10_cal = 16'b0000001111100110;
            15'd9665: log10_cal = 16'b0000001111100110;
            15'd9666: log10_cal = 16'b0000001111100110;
            15'd9667: log10_cal = 16'b0000001111100110;
            15'd9668: log10_cal = 16'b0000001111100110;
            15'd9669: log10_cal = 16'b0000001111100110;
            15'd9670: log10_cal = 16'b0000001111100110;
            15'd9671: log10_cal = 16'b0000001111100110;
            15'd9672: log10_cal = 16'b0000001111100110;
            15'd9673: log10_cal = 16'b0000001111100110;
            15'd9674: log10_cal = 16'b0000001111100110;
            15'd9675: log10_cal = 16'b0000001111100110;
            15'd9676: log10_cal = 16'b0000001111100110;
            15'd9677: log10_cal = 16'b0000001111100110;
            15'd9678: log10_cal = 16'b0000001111100110;
            15'd9679: log10_cal = 16'b0000001111100110;
            15'd9680: log10_cal = 16'b0000001111100110;
            15'd9681: log10_cal = 16'b0000001111100111;
            15'd9682: log10_cal = 16'b0000001111100111;
            15'd9683: log10_cal = 16'b0000001111100111;
            15'd9684: log10_cal = 16'b0000001111100111;
            15'd9685: log10_cal = 16'b0000001111100111;
            15'd9686: log10_cal = 16'b0000001111100111;
            15'd9687: log10_cal = 16'b0000001111100111;
            15'd9688: log10_cal = 16'b0000001111100111;
            15'd9689: log10_cal = 16'b0000001111100111;
            15'd9690: log10_cal = 16'b0000001111100111;
            15'd9691: log10_cal = 16'b0000001111100111;
            15'd9692: log10_cal = 16'b0000001111100111;
            15'd9693: log10_cal = 16'b0000001111100111;
            15'd9694: log10_cal = 16'b0000001111100111;
            15'd9695: log10_cal = 16'b0000001111100111;
            15'd9696: log10_cal = 16'b0000001111100111;
            15'd9697: log10_cal = 16'b0000001111100111;
            15'd9698: log10_cal = 16'b0000001111100111;
            15'd9699: log10_cal = 16'b0000001111100111;
            15'd9700: log10_cal = 16'b0000001111100111;
            15'd9701: log10_cal = 16'b0000001111100111;
            15'd9702: log10_cal = 16'b0000001111100111;
            15'd9703: log10_cal = 16'b0000001111101000;
            15'd9704: log10_cal = 16'b0000001111101000;
            15'd9705: log10_cal = 16'b0000001111101000;
            15'd9706: log10_cal = 16'b0000001111101000;
            15'd9707: log10_cal = 16'b0000001111101000;
            15'd9708: log10_cal = 16'b0000001111101000;
            15'd9709: log10_cal = 16'b0000001111101000;
            15'd9710: log10_cal = 16'b0000001111101000;
            15'd9711: log10_cal = 16'b0000001111101000;
            15'd9712: log10_cal = 16'b0000001111101000;
            15'd9713: log10_cal = 16'b0000001111101000;
            15'd9714: log10_cal = 16'b0000001111101000;
            15'd9715: log10_cal = 16'b0000001111101000;
            15'd9716: log10_cal = 16'b0000001111101000;
            15'd9717: log10_cal = 16'b0000001111101000;
            15'd9718: log10_cal = 16'b0000001111101000;
            15'd9719: log10_cal = 16'b0000001111101000;
            15'd9720: log10_cal = 16'b0000001111101000;
            15'd9721: log10_cal = 16'b0000001111101000;
            15'd9722: log10_cal = 16'b0000001111101000;
            15'd9723: log10_cal = 16'b0000001111101000;
            15'd9724: log10_cal = 16'b0000001111101001;
            15'd9725: log10_cal = 16'b0000001111101001;
            15'd9726: log10_cal = 16'b0000001111101001;
            15'd9727: log10_cal = 16'b0000001111101001;
            15'd9728: log10_cal = 16'b0000001111101001;
            15'd9729: log10_cal = 16'b0000001111101001;
            15'd9730: log10_cal = 16'b0000001111101001;
            15'd9731: log10_cal = 16'b0000001111101001;
            15'd9732: log10_cal = 16'b0000001111101001;
            15'd9733: log10_cal = 16'b0000001111101001;
            15'd9734: log10_cal = 16'b0000001111101001;
            15'd9735: log10_cal = 16'b0000001111101001;
            15'd9736: log10_cal = 16'b0000001111101001;
            15'd9737: log10_cal = 16'b0000001111101001;
            15'd9738: log10_cal = 16'b0000001111101001;
            15'd9739: log10_cal = 16'b0000001111101001;
            15'd9740: log10_cal = 16'b0000001111101001;
            15'd9741: log10_cal = 16'b0000001111101001;
            15'd9742: log10_cal = 16'b0000001111101001;
            15'd9743: log10_cal = 16'b0000001111101001;
            15'd9744: log10_cal = 16'b0000001111101001;
            15'd9745: log10_cal = 16'b0000001111101001;
            15'd9746: log10_cal = 16'b0000001111101010;
            15'd9747: log10_cal = 16'b0000001111101010;
            15'd9748: log10_cal = 16'b0000001111101010;
            15'd9749: log10_cal = 16'b0000001111101010;
            15'd9750: log10_cal = 16'b0000001111101010;
            15'd9751: log10_cal = 16'b0000001111101010;
            15'd9752: log10_cal = 16'b0000001111101010;
            15'd9753: log10_cal = 16'b0000001111101010;
            15'd9754: log10_cal = 16'b0000001111101010;
            15'd9755: log10_cal = 16'b0000001111101010;
            15'd9756: log10_cal = 16'b0000001111101010;
            15'd9757: log10_cal = 16'b0000001111101010;
            15'd9758: log10_cal = 16'b0000001111101010;
            15'd9759: log10_cal = 16'b0000001111101010;
            15'd9760: log10_cal = 16'b0000001111101010;
            15'd9761: log10_cal = 16'b0000001111101010;
            15'd9762: log10_cal = 16'b0000001111101010;
            15'd9763: log10_cal = 16'b0000001111101010;
            15'd9764: log10_cal = 16'b0000001111101010;
            15'd9765: log10_cal = 16'b0000001111101010;
            15'd9766: log10_cal = 16'b0000001111101010;
            15'd9767: log10_cal = 16'b0000001111101010;
            15'd9768: log10_cal = 16'b0000001111101011;
            15'd9769: log10_cal = 16'b0000001111101011;
            15'd9770: log10_cal = 16'b0000001111101011;
            15'd9771: log10_cal = 16'b0000001111101011;
            15'd9772: log10_cal = 16'b0000001111101011;
            15'd9773: log10_cal = 16'b0000001111101011;
            15'd9774: log10_cal = 16'b0000001111101011;
            15'd9775: log10_cal = 16'b0000001111101011;
            15'd9776: log10_cal = 16'b0000001111101011;
            15'd9777: log10_cal = 16'b0000001111101011;
            15'd9778: log10_cal = 16'b0000001111101011;
            15'd9779: log10_cal = 16'b0000001111101011;
            15'd9780: log10_cal = 16'b0000001111101011;
            15'd9781: log10_cal = 16'b0000001111101011;
            15'd9782: log10_cal = 16'b0000001111101011;
            15'd9783: log10_cal = 16'b0000001111101011;
            15'd9784: log10_cal = 16'b0000001111101011;
            15'd9785: log10_cal = 16'b0000001111101011;
            15'd9786: log10_cal = 16'b0000001111101011;
            15'd9787: log10_cal = 16'b0000001111101011;
            15'd9788: log10_cal = 16'b0000001111101011;
            15'd9789: log10_cal = 16'b0000001111101011;
            15'd9790: log10_cal = 16'b0000001111101100;
            15'd9791: log10_cal = 16'b0000001111101100;
            15'd9792: log10_cal = 16'b0000001111101100;
            15'd9793: log10_cal = 16'b0000001111101100;
            15'd9794: log10_cal = 16'b0000001111101100;
            15'd9795: log10_cal = 16'b0000001111101100;
            15'd9796: log10_cal = 16'b0000001111101100;
            15'd9797: log10_cal = 16'b0000001111101100;
            15'd9798: log10_cal = 16'b0000001111101100;
            15'd9799: log10_cal = 16'b0000001111101100;
            15'd9800: log10_cal = 16'b0000001111101100;
            15'd9801: log10_cal = 16'b0000001111101100;
            15'd9802: log10_cal = 16'b0000001111101100;
            15'd9803: log10_cal = 16'b0000001111101100;
            15'd9804: log10_cal = 16'b0000001111101100;
            15'd9805: log10_cal = 16'b0000001111101100;
            15'd9806: log10_cal = 16'b0000001111101100;
            15'd9807: log10_cal = 16'b0000001111101100;
            15'd9808: log10_cal = 16'b0000001111101100;
            15'd9809: log10_cal = 16'b0000001111101100;
            15'd9810: log10_cal = 16'b0000001111101100;
            15'd9811: log10_cal = 16'b0000001111101100;
            15'd9812: log10_cal = 16'b0000001111101101;
            15'd9813: log10_cal = 16'b0000001111101101;
            15'd9814: log10_cal = 16'b0000001111101101;
            15'd9815: log10_cal = 16'b0000001111101101;
            15'd9816: log10_cal = 16'b0000001111101101;
            15'd9817: log10_cal = 16'b0000001111101101;
            15'd9818: log10_cal = 16'b0000001111101101;
            15'd9819: log10_cal = 16'b0000001111101101;
            15'd9820: log10_cal = 16'b0000001111101101;
            15'd9821: log10_cal = 16'b0000001111101101;
            15'd9822: log10_cal = 16'b0000001111101101;
            15'd9823: log10_cal = 16'b0000001111101101;
            15'd9824: log10_cal = 16'b0000001111101101;
            15'd9825: log10_cal = 16'b0000001111101101;
            15'd9826: log10_cal = 16'b0000001111101101;
            15'd9827: log10_cal = 16'b0000001111101101;
            15'd9828: log10_cal = 16'b0000001111101101;
            15'd9829: log10_cal = 16'b0000001111101101;
            15'd9830: log10_cal = 16'b0000001111101101;
            15'd9831: log10_cal = 16'b0000001111101101;
            15'd9832: log10_cal = 16'b0000001111101101;
            15'd9833: log10_cal = 16'b0000001111101101;
            15'd9834: log10_cal = 16'b0000001111101110;
            15'd9835: log10_cal = 16'b0000001111101110;
            15'd9836: log10_cal = 16'b0000001111101110;
            15'd9837: log10_cal = 16'b0000001111101110;
            15'd9838: log10_cal = 16'b0000001111101110;
            15'd9839: log10_cal = 16'b0000001111101110;
            15'd9840: log10_cal = 16'b0000001111101110;
            15'd9841: log10_cal = 16'b0000001111101110;
            15'd9842: log10_cal = 16'b0000001111101110;
            15'd9843: log10_cal = 16'b0000001111101110;
            15'd9844: log10_cal = 16'b0000001111101110;
            15'd9845: log10_cal = 16'b0000001111101110;
            15'd9846: log10_cal = 16'b0000001111101110;
            15'd9847: log10_cal = 16'b0000001111101110;
            15'd9848: log10_cal = 16'b0000001111101110;
            15'd9849: log10_cal = 16'b0000001111101110;
            15'd9850: log10_cal = 16'b0000001111101110;
            15'd9851: log10_cal = 16'b0000001111101110;
            15'd9852: log10_cal = 16'b0000001111101110;
            15'd9853: log10_cal = 16'b0000001111101110;
            15'd9854: log10_cal = 16'b0000001111101110;
            15'd9855: log10_cal = 16'b0000001111101110;
            15'd9856: log10_cal = 16'b0000001111101111;
            15'd9857: log10_cal = 16'b0000001111101111;
            15'd9858: log10_cal = 16'b0000001111101111;
            15'd9859: log10_cal = 16'b0000001111101111;
            15'd9860: log10_cal = 16'b0000001111101111;
            15'd9861: log10_cal = 16'b0000001111101111;
            15'd9862: log10_cal = 16'b0000001111101111;
            15'd9863: log10_cal = 16'b0000001111101111;
            15'd9864: log10_cal = 16'b0000001111101111;
            15'd9865: log10_cal = 16'b0000001111101111;
            15'd9866: log10_cal = 16'b0000001111101111;
            15'd9867: log10_cal = 16'b0000001111101111;
            15'd9868: log10_cal = 16'b0000001111101111;
            15'd9869: log10_cal = 16'b0000001111101111;
            15'd9870: log10_cal = 16'b0000001111101111;
            15'd9871: log10_cal = 16'b0000001111101111;
            15'd9872: log10_cal = 16'b0000001111101111;
            15'd9873: log10_cal = 16'b0000001111101111;
            15'd9874: log10_cal = 16'b0000001111101111;
            15'd9875: log10_cal = 16'b0000001111101111;
            15'd9876: log10_cal = 16'b0000001111101111;
            15'd9877: log10_cal = 16'b0000001111101111;
            15'd9878: log10_cal = 16'b0000001111101111;
            15'd9879: log10_cal = 16'b0000001111110000;
            15'd9880: log10_cal = 16'b0000001111110000;
            15'd9881: log10_cal = 16'b0000001111110000;
            15'd9882: log10_cal = 16'b0000001111110000;
            15'd9883: log10_cal = 16'b0000001111110000;
            15'd9884: log10_cal = 16'b0000001111110000;
            15'd9885: log10_cal = 16'b0000001111110000;
            15'd9886: log10_cal = 16'b0000001111110000;
            15'd9887: log10_cal = 16'b0000001111110000;
            15'd9888: log10_cal = 16'b0000001111110000;
            15'd9889: log10_cal = 16'b0000001111110000;
            15'd9890: log10_cal = 16'b0000001111110000;
            15'd9891: log10_cal = 16'b0000001111110000;
            15'd9892: log10_cal = 16'b0000001111110000;
            15'd9893: log10_cal = 16'b0000001111110000;
            15'd9894: log10_cal = 16'b0000001111110000;
            15'd9895: log10_cal = 16'b0000001111110000;
            15'd9896: log10_cal = 16'b0000001111110000;
            15'd9897: log10_cal = 16'b0000001111110000;
            15'd9898: log10_cal = 16'b0000001111110000;
            15'd9899: log10_cal = 16'b0000001111110000;
            15'd9900: log10_cal = 16'b0000001111110000;
            15'd9901: log10_cal = 16'b0000001111110001;
            15'd9902: log10_cal = 16'b0000001111110001;
            15'd9903: log10_cal = 16'b0000001111110001;
            15'd9904: log10_cal = 16'b0000001111110001;
            15'd9905: log10_cal = 16'b0000001111110001;
            15'd9906: log10_cal = 16'b0000001111110001;
            15'd9907: log10_cal = 16'b0000001111110001;
            15'd9908: log10_cal = 16'b0000001111110001;
            15'd9909: log10_cal = 16'b0000001111110001;
            15'd9910: log10_cal = 16'b0000001111110001;
            15'd9911: log10_cal = 16'b0000001111110001;
            15'd9912: log10_cal = 16'b0000001111110001;
            15'd9913: log10_cal = 16'b0000001111110001;
            15'd9914: log10_cal = 16'b0000001111110001;
            15'd9915: log10_cal = 16'b0000001111110001;
            15'd9916: log10_cal = 16'b0000001111110001;
            15'd9917: log10_cal = 16'b0000001111110001;
            15'd9918: log10_cal = 16'b0000001111110001;
            15'd9919: log10_cal = 16'b0000001111110001;
            15'd9920: log10_cal = 16'b0000001111110001;
            15'd9921: log10_cal = 16'b0000001111110001;
            15'd9922: log10_cal = 16'b0000001111110001;
            15'd9923: log10_cal = 16'b0000001111110010;
            15'd9924: log10_cal = 16'b0000001111110010;
            15'd9925: log10_cal = 16'b0000001111110010;
            15'd9926: log10_cal = 16'b0000001111110010;
            15'd9927: log10_cal = 16'b0000001111110010;
            15'd9928: log10_cal = 16'b0000001111110010;
            15'd9929: log10_cal = 16'b0000001111110010;
            15'd9930: log10_cal = 16'b0000001111110010;
            15'd9931: log10_cal = 16'b0000001111110010;
            15'd9932: log10_cal = 16'b0000001111110010;
            15'd9933: log10_cal = 16'b0000001111110010;
            15'd9934: log10_cal = 16'b0000001111110010;
            15'd9935: log10_cal = 16'b0000001111110010;
            15'd9936: log10_cal = 16'b0000001111110010;
            15'd9937: log10_cal = 16'b0000001111110010;
            15'd9938: log10_cal = 16'b0000001111110010;
            15'd9939: log10_cal = 16'b0000001111110010;
            15'd9940: log10_cal = 16'b0000001111110010;
            15'd9941: log10_cal = 16'b0000001111110010;
            15'd9942: log10_cal = 16'b0000001111110010;
            15'd9943: log10_cal = 16'b0000001111110010;
            15'd9944: log10_cal = 16'b0000001111110010;
            15'd9945: log10_cal = 16'b0000001111110011;
            15'd9946: log10_cal = 16'b0000001111110011;
            15'd9947: log10_cal = 16'b0000001111110011;
            15'd9948: log10_cal = 16'b0000001111110011;
            15'd9949: log10_cal = 16'b0000001111110011;
            15'd9950: log10_cal = 16'b0000001111110011;
            15'd9951: log10_cal = 16'b0000001111110011;
            15'd9952: log10_cal = 16'b0000001111110011;
            15'd9953: log10_cal = 16'b0000001111110011;
            15'd9954: log10_cal = 16'b0000001111110011;
            15'd9955: log10_cal = 16'b0000001111110011;
            15'd9956: log10_cal = 16'b0000001111110011;
            15'd9957: log10_cal = 16'b0000001111110011;
            15'd9958: log10_cal = 16'b0000001111110011;
            15'd9959: log10_cal = 16'b0000001111110011;
            15'd9960: log10_cal = 16'b0000001111110011;
            15'd9961: log10_cal = 16'b0000001111110011;
            15'd9962: log10_cal = 16'b0000001111110011;
            15'd9963: log10_cal = 16'b0000001111110011;
            15'd9964: log10_cal = 16'b0000001111110011;
            15'd9965: log10_cal = 16'b0000001111110011;
            15'd9966: log10_cal = 16'b0000001111110011;
            15'd9967: log10_cal = 16'b0000001111110011;
            15'd9968: log10_cal = 16'b0000001111110100;
            15'd9969: log10_cal = 16'b0000001111110100;
            15'd9970: log10_cal = 16'b0000001111110100;
            15'd9971: log10_cal = 16'b0000001111110100;
            15'd9972: log10_cal = 16'b0000001111110100;
            15'd9973: log10_cal = 16'b0000001111110100;
            15'd9974: log10_cal = 16'b0000001111110100;
            15'd9975: log10_cal = 16'b0000001111110100;
            15'd9976: log10_cal = 16'b0000001111110100;
            15'd9977: log10_cal = 16'b0000001111110100;
            15'd9978: log10_cal = 16'b0000001111110100;
            15'd9979: log10_cal = 16'b0000001111110100;
            15'd9980: log10_cal = 16'b0000001111110100;
            15'd9981: log10_cal = 16'b0000001111110100;
            15'd9982: log10_cal = 16'b0000001111110100;
            15'd9983: log10_cal = 16'b0000001111110100;
            15'd9984: log10_cal = 16'b0000001111110100;
            15'd9985: log10_cal = 16'b0000001111110100;
            15'd9986: log10_cal = 16'b0000001111110100;
            15'd9987: log10_cal = 16'b0000001111110100;
            15'd9988: log10_cal = 16'b0000001111110100;
            15'd9989: log10_cal = 16'b0000001111110100;
            15'd9990: log10_cal = 16'b0000001111110101;
            15'd9991: log10_cal = 16'b0000001111110101;
            15'd9992: log10_cal = 16'b0000001111110101;
            15'd9993: log10_cal = 16'b0000001111110101;
            15'd9994: log10_cal = 16'b0000001111110101;
            15'd9995: log10_cal = 16'b0000001111110101;
            15'd9996: log10_cal = 16'b0000001111110101;
            15'd9997: log10_cal = 16'b0000001111110101;
            15'd9998: log10_cal = 16'b0000001111110101;
            15'd9999: log10_cal = 16'b0000001111110101;
            15'd10000: log10_cal = 16'b0000001111110101;
            15'd10001: log10_cal = 16'b0000001111110101;
            15'd10002: log10_cal = 16'b0000001111110101;
            15'd10003: log10_cal = 16'b0000001111110101;
            15'd10004: log10_cal = 16'b0000001111110101;
            15'd10005: log10_cal = 16'b0000001111110101;
            15'd10006: log10_cal = 16'b0000001111110101;
            15'd10007: log10_cal = 16'b0000001111110101;
            15'd10008: log10_cal = 16'b0000001111110101;
            15'd10009: log10_cal = 16'b0000001111110101;
            15'd10010: log10_cal = 16'b0000001111110101;
            15'd10011: log10_cal = 16'b0000001111110101;
            15'd10012: log10_cal = 16'b0000001111110101;
            15'd10013: log10_cal = 16'b0000001111110110;
            15'd10014: log10_cal = 16'b0000001111110110;
            15'd10015: log10_cal = 16'b0000001111110110;
            15'd10016: log10_cal = 16'b0000001111110110;
            15'd10017: log10_cal = 16'b0000001111110110;
            15'd10018: log10_cal = 16'b0000001111110110;
            15'd10019: log10_cal = 16'b0000001111110110;
            15'd10020: log10_cal = 16'b0000001111110110;
            15'd10021: log10_cal = 16'b0000001111110110;
            15'd10022: log10_cal = 16'b0000001111110110;
            15'd10023: log10_cal = 16'b0000001111110110;
            15'd10024: log10_cal = 16'b0000001111110110;
            15'd10025: log10_cal = 16'b0000001111110110;
            15'd10026: log10_cal = 16'b0000001111110110;
            15'd10027: log10_cal = 16'b0000001111110110;
            15'd10028: log10_cal = 16'b0000001111110110;
            15'd10029: log10_cal = 16'b0000001111110110;
            15'd10030: log10_cal = 16'b0000001111110110;
            15'd10031: log10_cal = 16'b0000001111110110;
            15'd10032: log10_cal = 16'b0000001111110110;
            15'd10033: log10_cal = 16'b0000001111110110;
            15'd10034: log10_cal = 16'b0000001111110110;
            15'd10035: log10_cal = 16'b0000001111110111;
            15'd10036: log10_cal = 16'b0000001111110111;
            15'd10037: log10_cal = 16'b0000001111110111;
            15'd10038: log10_cal = 16'b0000001111110111;
            15'd10039: log10_cal = 16'b0000001111110111;
            15'd10040: log10_cal = 16'b0000001111110111;
            15'd10041: log10_cal = 16'b0000001111110111;
            15'd10042: log10_cal = 16'b0000001111110111;
            15'd10043: log10_cal = 16'b0000001111110111;
            15'd10044: log10_cal = 16'b0000001111110111;
            15'd10045: log10_cal = 16'b0000001111110111;
            15'd10046: log10_cal = 16'b0000001111110111;
            15'd10047: log10_cal = 16'b0000001111110111;
            15'd10048: log10_cal = 16'b0000001111110111;
            15'd10049: log10_cal = 16'b0000001111110111;
            15'd10050: log10_cal = 16'b0000001111110111;
            15'd10051: log10_cal = 16'b0000001111110111;
            15'd10052: log10_cal = 16'b0000001111110111;
            15'd10053: log10_cal = 16'b0000001111110111;
            15'd10054: log10_cal = 16'b0000001111110111;
            15'd10055: log10_cal = 16'b0000001111110111;
            15'd10056: log10_cal = 16'b0000001111110111;
            15'd10057: log10_cal = 16'b0000001111110111;
            15'd10058: log10_cal = 16'b0000001111111000;
            15'd10059: log10_cal = 16'b0000001111111000;
            15'd10060: log10_cal = 16'b0000001111111000;
            15'd10061: log10_cal = 16'b0000001111111000;
            15'd10062: log10_cal = 16'b0000001111111000;
            15'd10063: log10_cal = 16'b0000001111111000;
            15'd10064: log10_cal = 16'b0000001111111000;
            15'd10065: log10_cal = 16'b0000001111111000;
            15'd10066: log10_cal = 16'b0000001111111000;
            15'd10067: log10_cal = 16'b0000001111111000;
            15'd10068: log10_cal = 16'b0000001111111000;
            15'd10069: log10_cal = 16'b0000001111111000;
            15'd10070: log10_cal = 16'b0000001111111000;
            15'd10071: log10_cal = 16'b0000001111111000;
            15'd10072: log10_cal = 16'b0000001111111000;
            15'd10073: log10_cal = 16'b0000001111111000;
            15'd10074: log10_cal = 16'b0000001111111000;
            15'd10075: log10_cal = 16'b0000001111111000;
            15'd10076: log10_cal = 16'b0000001111111000;
            15'd10077: log10_cal = 16'b0000001111111000;
            15'd10078: log10_cal = 16'b0000001111111000;
            15'd10079: log10_cal = 16'b0000001111111000;
            15'd10080: log10_cal = 16'b0000001111111000;
            15'd10081: log10_cal = 16'b0000001111111001;
            15'd10082: log10_cal = 16'b0000001111111001;
            15'd10083: log10_cal = 16'b0000001111111001;
            15'd10084: log10_cal = 16'b0000001111111001;
            15'd10085: log10_cal = 16'b0000001111111001;
            15'd10086: log10_cal = 16'b0000001111111001;
            15'd10087: log10_cal = 16'b0000001111111001;
            15'd10088: log10_cal = 16'b0000001111111001;
            15'd10089: log10_cal = 16'b0000001111111001;
            15'd10090: log10_cal = 16'b0000001111111001;
            15'd10091: log10_cal = 16'b0000001111111001;
            15'd10092: log10_cal = 16'b0000001111111001;
            15'd10093: log10_cal = 16'b0000001111111001;
            15'd10094: log10_cal = 16'b0000001111111001;
            15'd10095: log10_cal = 16'b0000001111111001;
            15'd10096: log10_cal = 16'b0000001111111001;
            15'd10097: log10_cal = 16'b0000001111111001;
            15'd10098: log10_cal = 16'b0000001111111001;
            15'd10099: log10_cal = 16'b0000001111111001;
            15'd10100: log10_cal = 16'b0000001111111001;
            15'd10101: log10_cal = 16'b0000001111111001;
            15'd10102: log10_cal = 16'b0000001111111001;
            15'd10103: log10_cal = 16'b0000001111111010;
            15'd10104: log10_cal = 16'b0000001111111010;
            15'd10105: log10_cal = 16'b0000001111111010;
            15'd10106: log10_cal = 16'b0000001111111010;
            15'd10107: log10_cal = 16'b0000001111111010;
            15'd10108: log10_cal = 16'b0000001111111010;
            15'd10109: log10_cal = 16'b0000001111111010;
            15'd10110: log10_cal = 16'b0000001111111010;
            15'd10111: log10_cal = 16'b0000001111111010;
            15'd10112: log10_cal = 16'b0000001111111010;
            15'd10113: log10_cal = 16'b0000001111111010;
            15'd10114: log10_cal = 16'b0000001111111010;
            15'd10115: log10_cal = 16'b0000001111111010;
            15'd10116: log10_cal = 16'b0000001111111010;
            15'd10117: log10_cal = 16'b0000001111111010;
            15'd10118: log10_cal = 16'b0000001111111010;
            15'd10119: log10_cal = 16'b0000001111111010;
            15'd10120: log10_cal = 16'b0000001111111010;
            15'd10121: log10_cal = 16'b0000001111111010;
            15'd10122: log10_cal = 16'b0000001111111010;
            15'd10123: log10_cal = 16'b0000001111111010;
            15'd10124: log10_cal = 16'b0000001111111010;
            15'd10125: log10_cal = 16'b0000001111111010;
            15'd10126: log10_cal = 16'b0000001111111011;
            15'd10127: log10_cal = 16'b0000001111111011;
            15'd10128: log10_cal = 16'b0000001111111011;
            15'd10129: log10_cal = 16'b0000001111111011;
            15'd10130: log10_cal = 16'b0000001111111011;
            15'd10131: log10_cal = 16'b0000001111111011;
            15'd10132: log10_cal = 16'b0000001111111011;
            15'd10133: log10_cal = 16'b0000001111111011;
            15'd10134: log10_cal = 16'b0000001111111011;
            15'd10135: log10_cal = 16'b0000001111111011;
            15'd10136: log10_cal = 16'b0000001111111011;
            15'd10137: log10_cal = 16'b0000001111111011;
            15'd10138: log10_cal = 16'b0000001111111011;
            15'd10139: log10_cal = 16'b0000001111111011;
            15'd10140: log10_cal = 16'b0000001111111011;
            15'd10141: log10_cal = 16'b0000001111111011;
            15'd10142: log10_cal = 16'b0000001111111011;
            15'd10143: log10_cal = 16'b0000001111111011;
            15'd10144: log10_cal = 16'b0000001111111011;
            15'd10145: log10_cal = 16'b0000001111111011;
            15'd10146: log10_cal = 16'b0000001111111011;
            15'd10147: log10_cal = 16'b0000001111111011;
            15'd10148: log10_cal = 16'b0000001111111011;
            15'd10149: log10_cal = 16'b0000001111111100;
            15'd10150: log10_cal = 16'b0000001111111100;
            15'd10151: log10_cal = 16'b0000001111111100;
            15'd10152: log10_cal = 16'b0000001111111100;
            15'd10153: log10_cal = 16'b0000001111111100;
            15'd10154: log10_cal = 16'b0000001111111100;
            15'd10155: log10_cal = 16'b0000001111111100;
            15'd10156: log10_cal = 16'b0000001111111100;
            15'd10157: log10_cal = 16'b0000001111111100;
            15'd10158: log10_cal = 16'b0000001111111100;
            15'd10159: log10_cal = 16'b0000001111111100;
            15'd10160: log10_cal = 16'b0000001111111100;
            15'd10161: log10_cal = 16'b0000001111111100;
            15'd10162: log10_cal = 16'b0000001111111100;
            15'd10163: log10_cal = 16'b0000001111111100;
            15'd10164: log10_cal = 16'b0000001111111100;
            15'd10165: log10_cal = 16'b0000001111111100;
            15'd10166: log10_cal = 16'b0000001111111100;
            15'd10167: log10_cal = 16'b0000001111111100;
            15'd10168: log10_cal = 16'b0000001111111100;
            15'd10169: log10_cal = 16'b0000001111111100;
            15'd10170: log10_cal = 16'b0000001111111100;
            15'd10171: log10_cal = 16'b0000001111111100;
            15'd10172: log10_cal = 16'b0000001111111101;
            15'd10173: log10_cal = 16'b0000001111111101;
            15'd10174: log10_cal = 16'b0000001111111101;
            15'd10175: log10_cal = 16'b0000001111111101;
            15'd10176: log10_cal = 16'b0000001111111101;
            15'd10177: log10_cal = 16'b0000001111111101;
            15'd10178: log10_cal = 16'b0000001111111101;
            15'd10179: log10_cal = 16'b0000001111111101;
            15'd10180: log10_cal = 16'b0000001111111101;
            15'd10181: log10_cal = 16'b0000001111111101;
            15'd10182: log10_cal = 16'b0000001111111101;
            15'd10183: log10_cal = 16'b0000001111111101;
            15'd10184: log10_cal = 16'b0000001111111101;
            15'd10185: log10_cal = 16'b0000001111111101;
            15'd10186: log10_cal = 16'b0000001111111101;
            15'd10187: log10_cal = 16'b0000001111111101;
            15'd10188: log10_cal = 16'b0000001111111101;
            15'd10189: log10_cal = 16'b0000001111111101;
            15'd10190: log10_cal = 16'b0000001111111101;
            15'd10191: log10_cal = 16'b0000001111111101;
            15'd10192: log10_cal = 16'b0000001111111101;
            15'd10193: log10_cal = 16'b0000001111111101;
            15'd10194: log10_cal = 16'b0000001111111101;
            15'd10195: log10_cal = 16'b0000001111111110;
            15'd10196: log10_cal = 16'b0000001111111110;
            15'd10197: log10_cal = 16'b0000001111111110;
            15'd10198: log10_cal = 16'b0000001111111110;
            15'd10199: log10_cal = 16'b0000001111111110;
            15'd10200: log10_cal = 16'b0000001111111110;
            15'd10201: log10_cal = 16'b0000001111111110;
            15'd10202: log10_cal = 16'b0000001111111110;
            15'd10203: log10_cal = 16'b0000001111111110;
            15'd10204: log10_cal = 16'b0000001111111110;
            15'd10205: log10_cal = 16'b0000001111111110;
            15'd10206: log10_cal = 16'b0000001111111110;
            15'd10207: log10_cal = 16'b0000001111111110;
            15'd10208: log10_cal = 16'b0000001111111110;
            15'd10209: log10_cal = 16'b0000001111111110;
            15'd10210: log10_cal = 16'b0000001111111110;
            15'd10211: log10_cal = 16'b0000001111111110;
            15'd10212: log10_cal = 16'b0000001111111110;
            15'd10213: log10_cal = 16'b0000001111111110;
            15'd10214: log10_cal = 16'b0000001111111110;
            15'd10215: log10_cal = 16'b0000001111111110;
            15'd10216: log10_cal = 16'b0000001111111110;
            15'd10217: log10_cal = 16'b0000001111111110;
            15'd10218: log10_cal = 16'b0000001111111111;
            15'd10219: log10_cal = 16'b0000001111111111;
            15'd10220: log10_cal = 16'b0000001111111111;
            15'd10221: log10_cal = 16'b0000001111111111;
            15'd10222: log10_cal = 16'b0000001111111111;
            15'd10223: log10_cal = 16'b0000001111111111;
            15'd10224: log10_cal = 16'b0000001111111111;
            15'd10225: log10_cal = 16'b0000001111111111;
            15'd10226: log10_cal = 16'b0000001111111111;
            15'd10227: log10_cal = 16'b0000001111111111;
            15'd10228: log10_cal = 16'b0000001111111111;
            15'd10229: log10_cal = 16'b0000001111111111;
            15'd10230: log10_cal = 16'b0000001111111111;
            15'd10231: log10_cal = 16'b0000001111111111;
            15'd10232: log10_cal = 16'b0000001111111111;
            15'd10233: log10_cal = 16'b0000001111111111;
            15'd10234: log10_cal = 16'b0000001111111111;
            15'd10235: log10_cal = 16'b0000001111111111;
            15'd10236: log10_cal = 16'b0000001111111111;
            15'd10237: log10_cal = 16'b0000001111111111;
            15'd10238: log10_cal = 16'b0000001111111111;
            15'd10239: log10_cal = 16'b0000001111111111;
            15'd10240: log10_cal = 16'b0000010000000000;
            15'd10241: log10_cal = 16'b0000010000000000;
            15'd10242: log10_cal = 16'b0000010000000000;
            15'd10243: log10_cal = 16'b0000010000000000;
            15'd10244: log10_cal = 16'b0000010000000000;
            15'd10245: log10_cal = 16'b0000010000000000;
            15'd10246: log10_cal = 16'b0000010000000000;
            15'd10247: log10_cal = 16'b0000010000000000;
            15'd10248: log10_cal = 16'b0000010000000000;
            15'd10249: log10_cal = 16'b0000010000000000;
            15'd10250: log10_cal = 16'b0000010000000000;
            15'd10251: log10_cal = 16'b0000010000000000;
            15'd10252: log10_cal = 16'b0000010000000000;
            15'd10253: log10_cal = 16'b0000010000000000;
            15'd10254: log10_cal = 16'b0000010000000000;
            15'd10255: log10_cal = 16'b0000010000000000;
            15'd10256: log10_cal = 16'b0000010000000000;
            15'd10257: log10_cal = 16'b0000010000000000;
            15'd10258: log10_cal = 16'b0000010000000000;
            15'd10259: log10_cal = 16'b0000010000000000;
            15'd10260: log10_cal = 16'b0000010000000000;
            15'd10261: log10_cal = 16'b0000010000000000;
            15'd10262: log10_cal = 16'b0000010000000000;
            15'd10263: log10_cal = 16'b0000010000000000;
            15'd10264: log10_cal = 16'b0000010000000001;
            15'd10265: log10_cal = 16'b0000010000000001;
            15'd10266: log10_cal = 16'b0000010000000001;
            15'd10267: log10_cal = 16'b0000010000000001;
            15'd10268: log10_cal = 16'b0000010000000001;
            15'd10269: log10_cal = 16'b0000010000000001;
            15'd10270: log10_cal = 16'b0000010000000001;
            15'd10271: log10_cal = 16'b0000010000000001;
            15'd10272: log10_cal = 16'b0000010000000001;
            15'd10273: log10_cal = 16'b0000010000000001;
            15'd10274: log10_cal = 16'b0000010000000001;
            15'd10275: log10_cal = 16'b0000010000000001;
            15'd10276: log10_cal = 16'b0000010000000001;
            15'd10277: log10_cal = 16'b0000010000000001;
            15'd10278: log10_cal = 16'b0000010000000001;
            15'd10279: log10_cal = 16'b0000010000000001;
            15'd10280: log10_cal = 16'b0000010000000001;
            15'd10281: log10_cal = 16'b0000010000000001;
            15'd10282: log10_cal = 16'b0000010000000001;
            15'd10283: log10_cal = 16'b0000010000000001;
            15'd10284: log10_cal = 16'b0000010000000001;
            15'd10285: log10_cal = 16'b0000010000000001;
            15'd10286: log10_cal = 16'b0000010000000001;
            15'd10287: log10_cal = 16'b0000010000000010;
            15'd10288: log10_cal = 16'b0000010000000010;
            15'd10289: log10_cal = 16'b0000010000000010;
            15'd10290: log10_cal = 16'b0000010000000010;
            15'd10291: log10_cal = 16'b0000010000000010;
            15'd10292: log10_cal = 16'b0000010000000010;
            15'd10293: log10_cal = 16'b0000010000000010;
            15'd10294: log10_cal = 16'b0000010000000010;
            15'd10295: log10_cal = 16'b0000010000000010;
            15'd10296: log10_cal = 16'b0000010000000010;
            15'd10297: log10_cal = 16'b0000010000000010;
            15'd10298: log10_cal = 16'b0000010000000010;
            15'd10299: log10_cal = 16'b0000010000000010;
            15'd10300: log10_cal = 16'b0000010000000010;
            15'd10301: log10_cal = 16'b0000010000000010;
            15'd10302: log10_cal = 16'b0000010000000010;
            15'd10303: log10_cal = 16'b0000010000000010;
            15'd10304: log10_cal = 16'b0000010000000010;
            15'd10305: log10_cal = 16'b0000010000000010;
            15'd10306: log10_cal = 16'b0000010000000010;
            15'd10307: log10_cal = 16'b0000010000000010;
            15'd10308: log10_cal = 16'b0000010000000010;
            15'd10309: log10_cal = 16'b0000010000000010;
            15'd10310: log10_cal = 16'b0000010000000011;
            15'd10311: log10_cal = 16'b0000010000000011;
            15'd10312: log10_cal = 16'b0000010000000011;
            15'd10313: log10_cal = 16'b0000010000000011;
            15'd10314: log10_cal = 16'b0000010000000011;
            15'd10315: log10_cal = 16'b0000010000000011;
            15'd10316: log10_cal = 16'b0000010000000011;
            15'd10317: log10_cal = 16'b0000010000000011;
            15'd10318: log10_cal = 16'b0000010000000011;
            15'd10319: log10_cal = 16'b0000010000000011;
            15'd10320: log10_cal = 16'b0000010000000011;
            15'd10321: log10_cal = 16'b0000010000000011;
            15'd10322: log10_cal = 16'b0000010000000011;
            15'd10323: log10_cal = 16'b0000010000000011;
            15'd10324: log10_cal = 16'b0000010000000011;
            15'd10325: log10_cal = 16'b0000010000000011;
            15'd10326: log10_cal = 16'b0000010000000011;
            15'd10327: log10_cal = 16'b0000010000000011;
            15'd10328: log10_cal = 16'b0000010000000011;
            15'd10329: log10_cal = 16'b0000010000000011;
            15'd10330: log10_cal = 16'b0000010000000011;
            15'd10331: log10_cal = 16'b0000010000000011;
            15'd10332: log10_cal = 16'b0000010000000011;
            15'd10333: log10_cal = 16'b0000010000000100;
            15'd10334: log10_cal = 16'b0000010000000100;
            15'd10335: log10_cal = 16'b0000010000000100;
            15'd10336: log10_cal = 16'b0000010000000100;
            15'd10337: log10_cal = 16'b0000010000000100;
            15'd10338: log10_cal = 16'b0000010000000100;
            15'd10339: log10_cal = 16'b0000010000000100;
            15'd10340: log10_cal = 16'b0000010000000100;
            15'd10341: log10_cal = 16'b0000010000000100;
            15'd10342: log10_cal = 16'b0000010000000100;
            15'd10343: log10_cal = 16'b0000010000000100;
            15'd10344: log10_cal = 16'b0000010000000100;
            15'd10345: log10_cal = 16'b0000010000000100;
            15'd10346: log10_cal = 16'b0000010000000100;
            15'd10347: log10_cal = 16'b0000010000000100;
            15'd10348: log10_cal = 16'b0000010000000100;
            15'd10349: log10_cal = 16'b0000010000000100;
            15'd10350: log10_cal = 16'b0000010000000100;
            15'd10351: log10_cal = 16'b0000010000000100;
            15'd10352: log10_cal = 16'b0000010000000100;
            15'd10353: log10_cal = 16'b0000010000000100;
            15'd10354: log10_cal = 16'b0000010000000100;
            15'd10355: log10_cal = 16'b0000010000000100;
            15'd10356: log10_cal = 16'b0000010000000101;
            15'd10357: log10_cal = 16'b0000010000000101;
            15'd10358: log10_cal = 16'b0000010000000101;
            15'd10359: log10_cal = 16'b0000010000000101;
            15'd10360: log10_cal = 16'b0000010000000101;
            15'd10361: log10_cal = 16'b0000010000000101;
            15'd10362: log10_cal = 16'b0000010000000101;
            15'd10363: log10_cal = 16'b0000010000000101;
            15'd10364: log10_cal = 16'b0000010000000101;
            15'd10365: log10_cal = 16'b0000010000000101;
            15'd10366: log10_cal = 16'b0000010000000101;
            15'd10367: log10_cal = 16'b0000010000000101;
            15'd10368: log10_cal = 16'b0000010000000101;
            15'd10369: log10_cal = 16'b0000010000000101;
            15'd10370: log10_cal = 16'b0000010000000101;
            15'd10371: log10_cal = 16'b0000010000000101;
            15'd10372: log10_cal = 16'b0000010000000101;
            15'd10373: log10_cal = 16'b0000010000000101;
            15'd10374: log10_cal = 16'b0000010000000101;
            15'd10375: log10_cal = 16'b0000010000000101;
            15'd10376: log10_cal = 16'b0000010000000101;
            15'd10377: log10_cal = 16'b0000010000000101;
            15'd10378: log10_cal = 16'b0000010000000101;
            15'd10379: log10_cal = 16'b0000010000000101;
            15'd10380: log10_cal = 16'b0000010000000110;
            15'd10381: log10_cal = 16'b0000010000000110;
            15'd10382: log10_cal = 16'b0000010000000110;
            15'd10383: log10_cal = 16'b0000010000000110;
            15'd10384: log10_cal = 16'b0000010000000110;
            15'd10385: log10_cal = 16'b0000010000000110;
            15'd10386: log10_cal = 16'b0000010000000110;
            15'd10387: log10_cal = 16'b0000010000000110;
            15'd10388: log10_cal = 16'b0000010000000110;
            15'd10389: log10_cal = 16'b0000010000000110;
            15'd10390: log10_cal = 16'b0000010000000110;
            15'd10391: log10_cal = 16'b0000010000000110;
            15'd10392: log10_cal = 16'b0000010000000110;
            15'd10393: log10_cal = 16'b0000010000000110;
            15'd10394: log10_cal = 16'b0000010000000110;
            15'd10395: log10_cal = 16'b0000010000000110;
            15'd10396: log10_cal = 16'b0000010000000110;
            15'd10397: log10_cal = 16'b0000010000000110;
            15'd10398: log10_cal = 16'b0000010000000110;
            15'd10399: log10_cal = 16'b0000010000000110;
            15'd10400: log10_cal = 16'b0000010000000110;
            15'd10401: log10_cal = 16'b0000010000000110;
            15'd10402: log10_cal = 16'b0000010000000110;
            15'd10403: log10_cal = 16'b0000010000000111;
            15'd10404: log10_cal = 16'b0000010000000111;
            15'd10405: log10_cal = 16'b0000010000000111;
            15'd10406: log10_cal = 16'b0000010000000111;
            15'd10407: log10_cal = 16'b0000010000000111;
            15'd10408: log10_cal = 16'b0000010000000111;
            15'd10409: log10_cal = 16'b0000010000000111;
            15'd10410: log10_cal = 16'b0000010000000111;
            15'd10411: log10_cal = 16'b0000010000000111;
            15'd10412: log10_cal = 16'b0000010000000111;
            15'd10413: log10_cal = 16'b0000010000000111;
            15'd10414: log10_cal = 16'b0000010000000111;
            15'd10415: log10_cal = 16'b0000010000000111;
            15'd10416: log10_cal = 16'b0000010000000111;
            15'd10417: log10_cal = 16'b0000010000000111;
            15'd10418: log10_cal = 16'b0000010000000111;
            15'd10419: log10_cal = 16'b0000010000000111;
            15'd10420: log10_cal = 16'b0000010000000111;
            15'd10421: log10_cal = 16'b0000010000000111;
            15'd10422: log10_cal = 16'b0000010000000111;
            15'd10423: log10_cal = 16'b0000010000000111;
            15'd10424: log10_cal = 16'b0000010000000111;
            15'd10425: log10_cal = 16'b0000010000000111;
            15'd10426: log10_cal = 16'b0000010000001000;
            15'd10427: log10_cal = 16'b0000010000001000;
            15'd10428: log10_cal = 16'b0000010000001000;
            15'd10429: log10_cal = 16'b0000010000001000;
            15'd10430: log10_cal = 16'b0000010000001000;
            15'd10431: log10_cal = 16'b0000010000001000;
            15'd10432: log10_cal = 16'b0000010000001000;
            15'd10433: log10_cal = 16'b0000010000001000;
            15'd10434: log10_cal = 16'b0000010000001000;
            15'd10435: log10_cal = 16'b0000010000001000;
            15'd10436: log10_cal = 16'b0000010000001000;
            15'd10437: log10_cal = 16'b0000010000001000;
            15'd10438: log10_cal = 16'b0000010000001000;
            15'd10439: log10_cal = 16'b0000010000001000;
            15'd10440: log10_cal = 16'b0000010000001000;
            15'd10441: log10_cal = 16'b0000010000001000;
            15'd10442: log10_cal = 16'b0000010000001000;
            15'd10443: log10_cal = 16'b0000010000001000;
            15'd10444: log10_cal = 16'b0000010000001000;
            15'd10445: log10_cal = 16'b0000010000001000;
            15'd10446: log10_cal = 16'b0000010000001000;
            15'd10447: log10_cal = 16'b0000010000001000;
            15'd10448: log10_cal = 16'b0000010000001000;
            15'd10449: log10_cal = 16'b0000010000001000;
            15'd10450: log10_cal = 16'b0000010000001001;
            15'd10451: log10_cal = 16'b0000010000001001;
            15'd10452: log10_cal = 16'b0000010000001001;
            15'd10453: log10_cal = 16'b0000010000001001;
            15'd10454: log10_cal = 16'b0000010000001001;
            15'd10455: log10_cal = 16'b0000010000001001;
            15'd10456: log10_cal = 16'b0000010000001001;
            15'd10457: log10_cal = 16'b0000010000001001;
            15'd10458: log10_cal = 16'b0000010000001001;
            15'd10459: log10_cal = 16'b0000010000001001;
            15'd10460: log10_cal = 16'b0000010000001001;
            15'd10461: log10_cal = 16'b0000010000001001;
            15'd10462: log10_cal = 16'b0000010000001001;
            15'd10463: log10_cal = 16'b0000010000001001;
            15'd10464: log10_cal = 16'b0000010000001001;
            15'd10465: log10_cal = 16'b0000010000001001;
            15'd10466: log10_cal = 16'b0000010000001001;
            15'd10467: log10_cal = 16'b0000010000001001;
            15'd10468: log10_cal = 16'b0000010000001001;
            15'd10469: log10_cal = 16'b0000010000001001;
            15'd10470: log10_cal = 16'b0000010000001001;
            15'd10471: log10_cal = 16'b0000010000001001;
            15'd10472: log10_cal = 16'b0000010000001001;
            15'd10473: log10_cal = 16'b0000010000001010;
            15'd10474: log10_cal = 16'b0000010000001010;
            15'd10475: log10_cal = 16'b0000010000001010;
            15'd10476: log10_cal = 16'b0000010000001010;
            15'd10477: log10_cal = 16'b0000010000001010;
            15'd10478: log10_cal = 16'b0000010000001010;
            15'd10479: log10_cal = 16'b0000010000001010;
            15'd10480: log10_cal = 16'b0000010000001010;
            15'd10481: log10_cal = 16'b0000010000001010;
            15'd10482: log10_cal = 16'b0000010000001010;
            15'd10483: log10_cal = 16'b0000010000001010;
            15'd10484: log10_cal = 16'b0000010000001010;
            15'd10485: log10_cal = 16'b0000010000001010;
            15'd10486: log10_cal = 16'b0000010000001010;
            15'd10487: log10_cal = 16'b0000010000001010;
            15'd10488: log10_cal = 16'b0000010000001010;
            15'd10489: log10_cal = 16'b0000010000001010;
            15'd10490: log10_cal = 16'b0000010000001010;
            15'd10491: log10_cal = 16'b0000010000001010;
            15'd10492: log10_cal = 16'b0000010000001010;
            15'd10493: log10_cal = 16'b0000010000001010;
            15'd10494: log10_cal = 16'b0000010000001010;
            15'd10495: log10_cal = 16'b0000010000001010;
            15'd10496: log10_cal = 16'b0000010000001010;
            15'd10497: log10_cal = 16'b0000010000001011;
            15'd10498: log10_cal = 16'b0000010000001011;
            15'd10499: log10_cal = 16'b0000010000001011;
            15'd10500: log10_cal = 16'b0000010000001011;
            15'd10501: log10_cal = 16'b0000010000001011;
            15'd10502: log10_cal = 16'b0000010000001011;
            15'd10503: log10_cal = 16'b0000010000001011;
            15'd10504: log10_cal = 16'b0000010000001011;
            15'd10505: log10_cal = 16'b0000010000001011;
            15'd10506: log10_cal = 16'b0000010000001011;
            15'd10507: log10_cal = 16'b0000010000001011;
            15'd10508: log10_cal = 16'b0000010000001011;
            15'd10509: log10_cal = 16'b0000010000001011;
            15'd10510: log10_cal = 16'b0000010000001011;
            15'd10511: log10_cal = 16'b0000010000001011;
            15'd10512: log10_cal = 16'b0000010000001011;
            15'd10513: log10_cal = 16'b0000010000001011;
            15'd10514: log10_cal = 16'b0000010000001011;
            15'd10515: log10_cal = 16'b0000010000001011;
            15'd10516: log10_cal = 16'b0000010000001011;
            15'd10517: log10_cal = 16'b0000010000001011;
            15'd10518: log10_cal = 16'b0000010000001011;
            15'd10519: log10_cal = 16'b0000010000001011;
            15'd10520: log10_cal = 16'b0000010000001011;
            15'd10521: log10_cal = 16'b0000010000001100;
            15'd10522: log10_cal = 16'b0000010000001100;
            15'd10523: log10_cal = 16'b0000010000001100;
            15'd10524: log10_cal = 16'b0000010000001100;
            15'd10525: log10_cal = 16'b0000010000001100;
            15'd10526: log10_cal = 16'b0000010000001100;
            15'd10527: log10_cal = 16'b0000010000001100;
            15'd10528: log10_cal = 16'b0000010000001100;
            15'd10529: log10_cal = 16'b0000010000001100;
            15'd10530: log10_cal = 16'b0000010000001100;
            15'd10531: log10_cal = 16'b0000010000001100;
            15'd10532: log10_cal = 16'b0000010000001100;
            15'd10533: log10_cal = 16'b0000010000001100;
            15'd10534: log10_cal = 16'b0000010000001100;
            15'd10535: log10_cal = 16'b0000010000001100;
            15'd10536: log10_cal = 16'b0000010000001100;
            15'd10537: log10_cal = 16'b0000010000001100;
            15'd10538: log10_cal = 16'b0000010000001100;
            15'd10539: log10_cal = 16'b0000010000001100;
            15'd10540: log10_cal = 16'b0000010000001100;
            15'd10541: log10_cal = 16'b0000010000001100;
            15'd10542: log10_cal = 16'b0000010000001100;
            15'd10543: log10_cal = 16'b0000010000001100;
            15'd10544: log10_cal = 16'b0000010000001101;
            15'd10545: log10_cal = 16'b0000010000001101;
            15'd10546: log10_cal = 16'b0000010000001101;
            15'd10547: log10_cal = 16'b0000010000001101;
            15'd10548: log10_cal = 16'b0000010000001101;
            15'd10549: log10_cal = 16'b0000010000001101;
            15'd10550: log10_cal = 16'b0000010000001101;
            15'd10551: log10_cal = 16'b0000010000001101;
            15'd10552: log10_cal = 16'b0000010000001101;
            15'd10553: log10_cal = 16'b0000010000001101;
            15'd10554: log10_cal = 16'b0000010000001101;
            15'd10555: log10_cal = 16'b0000010000001101;
            15'd10556: log10_cal = 16'b0000010000001101;
            15'd10557: log10_cal = 16'b0000010000001101;
            15'd10558: log10_cal = 16'b0000010000001101;
            15'd10559: log10_cal = 16'b0000010000001101;
            15'd10560: log10_cal = 16'b0000010000001101;
            15'd10561: log10_cal = 16'b0000010000001101;
            15'd10562: log10_cal = 16'b0000010000001101;
            15'd10563: log10_cal = 16'b0000010000001101;
            15'd10564: log10_cal = 16'b0000010000001101;
            15'd10565: log10_cal = 16'b0000010000001101;
            15'd10566: log10_cal = 16'b0000010000001101;
            15'd10567: log10_cal = 16'b0000010000001101;
            15'd10568: log10_cal = 16'b0000010000001110;
            15'd10569: log10_cal = 16'b0000010000001110;
            15'd10570: log10_cal = 16'b0000010000001110;
            15'd10571: log10_cal = 16'b0000010000001110;
            15'd10572: log10_cal = 16'b0000010000001110;
            15'd10573: log10_cal = 16'b0000010000001110;
            15'd10574: log10_cal = 16'b0000010000001110;
            15'd10575: log10_cal = 16'b0000010000001110;
            15'd10576: log10_cal = 16'b0000010000001110;
            15'd10577: log10_cal = 16'b0000010000001110;
            15'd10578: log10_cal = 16'b0000010000001110;
            15'd10579: log10_cal = 16'b0000010000001110;
            15'd10580: log10_cal = 16'b0000010000001110;
            15'd10581: log10_cal = 16'b0000010000001110;
            15'd10582: log10_cal = 16'b0000010000001110;
            15'd10583: log10_cal = 16'b0000010000001110;
            15'd10584: log10_cal = 16'b0000010000001110;
            15'd10585: log10_cal = 16'b0000010000001110;
            15'd10586: log10_cal = 16'b0000010000001110;
            15'd10587: log10_cal = 16'b0000010000001110;
            15'd10588: log10_cal = 16'b0000010000001110;
            15'd10589: log10_cal = 16'b0000010000001110;
            15'd10590: log10_cal = 16'b0000010000001110;
            15'd10591: log10_cal = 16'b0000010000001110;
            15'd10592: log10_cal = 16'b0000010000001111;
            15'd10593: log10_cal = 16'b0000010000001111;
            15'd10594: log10_cal = 16'b0000010000001111;
            15'd10595: log10_cal = 16'b0000010000001111;
            15'd10596: log10_cal = 16'b0000010000001111;
            15'd10597: log10_cal = 16'b0000010000001111;
            15'd10598: log10_cal = 16'b0000010000001111;
            15'd10599: log10_cal = 16'b0000010000001111;
            15'd10600: log10_cal = 16'b0000010000001111;
            15'd10601: log10_cal = 16'b0000010000001111;
            15'd10602: log10_cal = 16'b0000010000001111;
            15'd10603: log10_cal = 16'b0000010000001111;
            15'd10604: log10_cal = 16'b0000010000001111;
            15'd10605: log10_cal = 16'b0000010000001111;
            15'd10606: log10_cal = 16'b0000010000001111;
            15'd10607: log10_cal = 16'b0000010000001111;
            15'd10608: log10_cal = 16'b0000010000001111;
            15'd10609: log10_cal = 16'b0000010000001111;
            15'd10610: log10_cal = 16'b0000010000001111;
            15'd10611: log10_cal = 16'b0000010000001111;
            15'd10612: log10_cal = 16'b0000010000001111;
            15'd10613: log10_cal = 16'b0000010000001111;
            15'd10614: log10_cal = 16'b0000010000001111;
            15'd10615: log10_cal = 16'b0000010000001111;
            15'd10616: log10_cal = 16'b0000010000010000;
            15'd10617: log10_cal = 16'b0000010000010000;
            15'd10618: log10_cal = 16'b0000010000010000;
            15'd10619: log10_cal = 16'b0000010000010000;
            15'd10620: log10_cal = 16'b0000010000010000;
            15'd10621: log10_cal = 16'b0000010000010000;
            15'd10622: log10_cal = 16'b0000010000010000;
            15'd10623: log10_cal = 16'b0000010000010000;
            15'd10624: log10_cal = 16'b0000010000010000;
            15'd10625: log10_cal = 16'b0000010000010000;
            15'd10626: log10_cal = 16'b0000010000010000;
            15'd10627: log10_cal = 16'b0000010000010000;
            15'd10628: log10_cal = 16'b0000010000010000;
            15'd10629: log10_cal = 16'b0000010000010000;
            15'd10630: log10_cal = 16'b0000010000010000;
            15'd10631: log10_cal = 16'b0000010000010000;
            15'd10632: log10_cal = 16'b0000010000010000;
            15'd10633: log10_cal = 16'b0000010000010000;
            15'd10634: log10_cal = 16'b0000010000010000;
            15'd10635: log10_cal = 16'b0000010000010000;
            15'd10636: log10_cal = 16'b0000010000010000;
            15'd10637: log10_cal = 16'b0000010000010000;
            15'd10638: log10_cal = 16'b0000010000010000;
            15'd10639: log10_cal = 16'b0000010000010000;
            15'd10640: log10_cal = 16'b0000010000010001;
            15'd10641: log10_cal = 16'b0000010000010001;
            15'd10642: log10_cal = 16'b0000010000010001;
            15'd10643: log10_cal = 16'b0000010000010001;
            15'd10644: log10_cal = 16'b0000010000010001;
            15'd10645: log10_cal = 16'b0000010000010001;
            15'd10646: log10_cal = 16'b0000010000010001;
            15'd10647: log10_cal = 16'b0000010000010001;
            15'd10648: log10_cal = 16'b0000010000010001;
            15'd10649: log10_cal = 16'b0000010000010001;
            15'd10650: log10_cal = 16'b0000010000010001;
            15'd10651: log10_cal = 16'b0000010000010001;
            15'd10652: log10_cal = 16'b0000010000010001;
            15'd10653: log10_cal = 16'b0000010000010001;
            15'd10654: log10_cal = 16'b0000010000010001;
            15'd10655: log10_cal = 16'b0000010000010001;
            15'd10656: log10_cal = 16'b0000010000010001;
            15'd10657: log10_cal = 16'b0000010000010001;
            15'd10658: log10_cal = 16'b0000010000010001;
            15'd10659: log10_cal = 16'b0000010000010001;
            15'd10660: log10_cal = 16'b0000010000010001;
            15'd10661: log10_cal = 16'b0000010000010001;
            15'd10662: log10_cal = 16'b0000010000010001;
            15'd10663: log10_cal = 16'b0000010000010010;
            15'd10664: log10_cal = 16'b0000010000010010;
            15'd10665: log10_cal = 16'b0000010000010010;
            15'd10666: log10_cal = 16'b0000010000010010;
            15'd10667: log10_cal = 16'b0000010000010010;
            15'd10668: log10_cal = 16'b0000010000010010;
            15'd10669: log10_cal = 16'b0000010000010010;
            15'd10670: log10_cal = 16'b0000010000010010;
            15'd10671: log10_cal = 16'b0000010000010010;
            15'd10672: log10_cal = 16'b0000010000010010;
            15'd10673: log10_cal = 16'b0000010000010010;
            15'd10674: log10_cal = 16'b0000010000010010;
            15'd10675: log10_cal = 16'b0000010000010010;
            15'd10676: log10_cal = 16'b0000010000010010;
            15'd10677: log10_cal = 16'b0000010000010010;
            15'd10678: log10_cal = 16'b0000010000010010;
            15'd10679: log10_cal = 16'b0000010000010010;
            15'd10680: log10_cal = 16'b0000010000010010;
            15'd10681: log10_cal = 16'b0000010000010010;
            15'd10682: log10_cal = 16'b0000010000010010;
            15'd10683: log10_cal = 16'b0000010000010010;
            15'd10684: log10_cal = 16'b0000010000010010;
            15'd10685: log10_cal = 16'b0000010000010010;
            15'd10686: log10_cal = 16'b0000010000010010;
            15'd10687: log10_cal = 16'b0000010000010011;
            15'd10688: log10_cal = 16'b0000010000010011;
            15'd10689: log10_cal = 16'b0000010000010011;
            15'd10690: log10_cal = 16'b0000010000010011;
            15'd10691: log10_cal = 16'b0000010000010011;
            15'd10692: log10_cal = 16'b0000010000010011;
            15'd10693: log10_cal = 16'b0000010000010011;
            15'd10694: log10_cal = 16'b0000010000010011;
            15'd10695: log10_cal = 16'b0000010000010011;
            15'd10696: log10_cal = 16'b0000010000010011;
            15'd10697: log10_cal = 16'b0000010000010011;
            15'd10698: log10_cal = 16'b0000010000010011;
            15'd10699: log10_cal = 16'b0000010000010011;
            15'd10700: log10_cal = 16'b0000010000010011;
            15'd10701: log10_cal = 16'b0000010000010011;
            15'd10702: log10_cal = 16'b0000010000010011;
            15'd10703: log10_cal = 16'b0000010000010011;
            15'd10704: log10_cal = 16'b0000010000010011;
            15'd10705: log10_cal = 16'b0000010000010011;
            15'd10706: log10_cal = 16'b0000010000010011;
            15'd10707: log10_cal = 16'b0000010000010011;
            15'd10708: log10_cal = 16'b0000010000010011;
            15'd10709: log10_cal = 16'b0000010000010011;
            15'd10710: log10_cal = 16'b0000010000010011;
            15'd10711: log10_cal = 16'b0000010000010011;
            15'd10712: log10_cal = 16'b0000010000010100;
            15'd10713: log10_cal = 16'b0000010000010100;
            15'd10714: log10_cal = 16'b0000010000010100;
            15'd10715: log10_cal = 16'b0000010000010100;
            15'd10716: log10_cal = 16'b0000010000010100;
            15'd10717: log10_cal = 16'b0000010000010100;
            15'd10718: log10_cal = 16'b0000010000010100;
            15'd10719: log10_cal = 16'b0000010000010100;
            15'd10720: log10_cal = 16'b0000010000010100;
            15'd10721: log10_cal = 16'b0000010000010100;
            15'd10722: log10_cal = 16'b0000010000010100;
            15'd10723: log10_cal = 16'b0000010000010100;
            15'd10724: log10_cal = 16'b0000010000010100;
            15'd10725: log10_cal = 16'b0000010000010100;
            15'd10726: log10_cal = 16'b0000010000010100;
            15'd10727: log10_cal = 16'b0000010000010100;
            15'd10728: log10_cal = 16'b0000010000010100;
            15'd10729: log10_cal = 16'b0000010000010100;
            15'd10730: log10_cal = 16'b0000010000010100;
            15'd10731: log10_cal = 16'b0000010000010100;
            15'd10732: log10_cal = 16'b0000010000010100;
            15'd10733: log10_cal = 16'b0000010000010100;
            15'd10734: log10_cal = 16'b0000010000010100;
            15'd10735: log10_cal = 16'b0000010000010100;
            15'd10736: log10_cal = 16'b0000010000010101;
            15'd10737: log10_cal = 16'b0000010000010101;
            15'd10738: log10_cal = 16'b0000010000010101;
            15'd10739: log10_cal = 16'b0000010000010101;
            15'd10740: log10_cal = 16'b0000010000010101;
            15'd10741: log10_cal = 16'b0000010000010101;
            15'd10742: log10_cal = 16'b0000010000010101;
            15'd10743: log10_cal = 16'b0000010000010101;
            15'd10744: log10_cal = 16'b0000010000010101;
            15'd10745: log10_cal = 16'b0000010000010101;
            15'd10746: log10_cal = 16'b0000010000010101;
            15'd10747: log10_cal = 16'b0000010000010101;
            15'd10748: log10_cal = 16'b0000010000010101;
            15'd10749: log10_cal = 16'b0000010000010101;
            15'd10750: log10_cal = 16'b0000010000010101;
            15'd10751: log10_cal = 16'b0000010000010101;
            15'd10752: log10_cal = 16'b0000010000010101;
            15'd10753: log10_cal = 16'b0000010000010101;
            15'd10754: log10_cal = 16'b0000010000010101;
            15'd10755: log10_cal = 16'b0000010000010101;
            15'd10756: log10_cal = 16'b0000010000010101;
            15'd10757: log10_cal = 16'b0000010000010101;
            15'd10758: log10_cal = 16'b0000010000010101;
            15'd10759: log10_cal = 16'b0000010000010101;
            15'd10760: log10_cal = 16'b0000010000010110;
            15'd10761: log10_cal = 16'b0000010000010110;
            15'd10762: log10_cal = 16'b0000010000010110;
            15'd10763: log10_cal = 16'b0000010000010110;
            15'd10764: log10_cal = 16'b0000010000010110;
            15'd10765: log10_cal = 16'b0000010000010110;
            15'd10766: log10_cal = 16'b0000010000010110;
            15'd10767: log10_cal = 16'b0000010000010110;
            15'd10768: log10_cal = 16'b0000010000010110;
            15'd10769: log10_cal = 16'b0000010000010110;
            15'd10770: log10_cal = 16'b0000010000010110;
            15'd10771: log10_cal = 16'b0000010000010110;
            15'd10772: log10_cal = 16'b0000010000010110;
            15'd10773: log10_cal = 16'b0000010000010110;
            15'd10774: log10_cal = 16'b0000010000010110;
            15'd10775: log10_cal = 16'b0000010000010110;
            15'd10776: log10_cal = 16'b0000010000010110;
            15'd10777: log10_cal = 16'b0000010000010110;
            15'd10778: log10_cal = 16'b0000010000010110;
            15'd10779: log10_cal = 16'b0000010000010110;
            15'd10780: log10_cal = 16'b0000010000010110;
            15'd10781: log10_cal = 16'b0000010000010110;
            15'd10782: log10_cal = 16'b0000010000010110;
            15'd10783: log10_cal = 16'b0000010000010110;
            15'd10784: log10_cal = 16'b0000010000010111;
            15'd10785: log10_cal = 16'b0000010000010111;
            15'd10786: log10_cal = 16'b0000010000010111;
            15'd10787: log10_cal = 16'b0000010000010111;
            15'd10788: log10_cal = 16'b0000010000010111;
            15'd10789: log10_cal = 16'b0000010000010111;
            15'd10790: log10_cal = 16'b0000010000010111;
            15'd10791: log10_cal = 16'b0000010000010111;
            15'd10792: log10_cal = 16'b0000010000010111;
            15'd10793: log10_cal = 16'b0000010000010111;
            15'd10794: log10_cal = 16'b0000010000010111;
            15'd10795: log10_cal = 16'b0000010000010111;
            15'd10796: log10_cal = 16'b0000010000010111;
            15'd10797: log10_cal = 16'b0000010000010111;
            15'd10798: log10_cal = 16'b0000010000010111;
            15'd10799: log10_cal = 16'b0000010000010111;
            15'd10800: log10_cal = 16'b0000010000010111;
            15'd10801: log10_cal = 16'b0000010000010111;
            15'd10802: log10_cal = 16'b0000010000010111;
            15'd10803: log10_cal = 16'b0000010000010111;
            15'd10804: log10_cal = 16'b0000010000010111;
            15'd10805: log10_cal = 16'b0000010000010111;
            15'd10806: log10_cal = 16'b0000010000010111;
            15'd10807: log10_cal = 16'b0000010000010111;
            15'd10808: log10_cal = 16'b0000010000011000;
            15'd10809: log10_cal = 16'b0000010000011000;
            15'd10810: log10_cal = 16'b0000010000011000;
            15'd10811: log10_cal = 16'b0000010000011000;
            15'd10812: log10_cal = 16'b0000010000011000;
            15'd10813: log10_cal = 16'b0000010000011000;
            15'd10814: log10_cal = 16'b0000010000011000;
            15'd10815: log10_cal = 16'b0000010000011000;
            15'd10816: log10_cal = 16'b0000010000011000;
            15'd10817: log10_cal = 16'b0000010000011000;
            15'd10818: log10_cal = 16'b0000010000011000;
            15'd10819: log10_cal = 16'b0000010000011000;
            15'd10820: log10_cal = 16'b0000010000011000;
            15'd10821: log10_cal = 16'b0000010000011000;
            15'd10822: log10_cal = 16'b0000010000011000;
            15'd10823: log10_cal = 16'b0000010000011000;
            15'd10824: log10_cal = 16'b0000010000011000;
            15'd10825: log10_cal = 16'b0000010000011000;
            15'd10826: log10_cal = 16'b0000010000011000;
            15'd10827: log10_cal = 16'b0000010000011000;
            15'd10828: log10_cal = 16'b0000010000011000;
            15'd10829: log10_cal = 16'b0000010000011000;
            15'd10830: log10_cal = 16'b0000010000011000;
            15'd10831: log10_cal = 16'b0000010000011000;
            15'd10832: log10_cal = 16'b0000010000011000;
            15'd10833: log10_cal = 16'b0000010000011001;
            15'd10834: log10_cal = 16'b0000010000011001;
            15'd10835: log10_cal = 16'b0000010000011001;
            15'd10836: log10_cal = 16'b0000010000011001;
            15'd10837: log10_cal = 16'b0000010000011001;
            15'd10838: log10_cal = 16'b0000010000011001;
            15'd10839: log10_cal = 16'b0000010000011001;
            15'd10840: log10_cal = 16'b0000010000011001;
            15'd10841: log10_cal = 16'b0000010000011001;
            15'd10842: log10_cal = 16'b0000010000011001;
            15'd10843: log10_cal = 16'b0000010000011001;
            15'd10844: log10_cal = 16'b0000010000011001;
            15'd10845: log10_cal = 16'b0000010000011001;
            15'd10846: log10_cal = 16'b0000010000011001;
            15'd10847: log10_cal = 16'b0000010000011001;
            15'd10848: log10_cal = 16'b0000010000011001;
            15'd10849: log10_cal = 16'b0000010000011001;
            15'd10850: log10_cal = 16'b0000010000011001;
            15'd10851: log10_cal = 16'b0000010000011001;
            15'd10852: log10_cal = 16'b0000010000011001;
            15'd10853: log10_cal = 16'b0000010000011001;
            15'd10854: log10_cal = 16'b0000010000011001;
            15'd10855: log10_cal = 16'b0000010000011001;
            15'd10856: log10_cal = 16'b0000010000011001;
            15'd10857: log10_cal = 16'b0000010000011010;
            15'd10858: log10_cal = 16'b0000010000011010;
            15'd10859: log10_cal = 16'b0000010000011010;
            15'd10860: log10_cal = 16'b0000010000011010;
            15'd10861: log10_cal = 16'b0000010000011010;
            15'd10862: log10_cal = 16'b0000010000011010;
            15'd10863: log10_cal = 16'b0000010000011010;
            15'd10864: log10_cal = 16'b0000010000011010;
            15'd10865: log10_cal = 16'b0000010000011010;
            15'd10866: log10_cal = 16'b0000010000011010;
            15'd10867: log10_cal = 16'b0000010000011010;
            15'd10868: log10_cal = 16'b0000010000011010;
            15'd10869: log10_cal = 16'b0000010000011010;
            15'd10870: log10_cal = 16'b0000010000011010;
            15'd10871: log10_cal = 16'b0000010000011010;
            15'd10872: log10_cal = 16'b0000010000011010;
            15'd10873: log10_cal = 16'b0000010000011010;
            15'd10874: log10_cal = 16'b0000010000011010;
            15'd10875: log10_cal = 16'b0000010000011010;
            15'd10876: log10_cal = 16'b0000010000011010;
            15'd10877: log10_cal = 16'b0000010000011010;
            15'd10878: log10_cal = 16'b0000010000011010;
            15'd10879: log10_cal = 16'b0000010000011010;
            15'd10880: log10_cal = 16'b0000010000011010;
            15'd10881: log10_cal = 16'b0000010000011011;
            15'd10882: log10_cal = 16'b0000010000011011;
            15'd10883: log10_cal = 16'b0000010000011011;
            15'd10884: log10_cal = 16'b0000010000011011;
            15'd10885: log10_cal = 16'b0000010000011011;
            15'd10886: log10_cal = 16'b0000010000011011;
            15'd10887: log10_cal = 16'b0000010000011011;
            15'd10888: log10_cal = 16'b0000010000011011;
            15'd10889: log10_cal = 16'b0000010000011011;
            15'd10890: log10_cal = 16'b0000010000011011;
            15'd10891: log10_cal = 16'b0000010000011011;
            15'd10892: log10_cal = 16'b0000010000011011;
            15'd10893: log10_cal = 16'b0000010000011011;
            15'd10894: log10_cal = 16'b0000010000011011;
            15'd10895: log10_cal = 16'b0000010000011011;
            15'd10896: log10_cal = 16'b0000010000011011;
            15'd10897: log10_cal = 16'b0000010000011011;
            15'd10898: log10_cal = 16'b0000010000011011;
            15'd10899: log10_cal = 16'b0000010000011011;
            15'd10900: log10_cal = 16'b0000010000011011;
            15'd10901: log10_cal = 16'b0000010000011011;
            15'd10902: log10_cal = 16'b0000010000011011;
            15'd10903: log10_cal = 16'b0000010000011011;
            15'd10904: log10_cal = 16'b0000010000011011;
            15'd10905: log10_cal = 16'b0000010000011011;
            15'd10906: log10_cal = 16'b0000010000011100;
            15'd10907: log10_cal = 16'b0000010000011100;
            15'd10908: log10_cal = 16'b0000010000011100;
            15'd10909: log10_cal = 16'b0000010000011100;
            15'd10910: log10_cal = 16'b0000010000011100;
            15'd10911: log10_cal = 16'b0000010000011100;
            15'd10912: log10_cal = 16'b0000010000011100;
            15'd10913: log10_cal = 16'b0000010000011100;
            15'd10914: log10_cal = 16'b0000010000011100;
            15'd10915: log10_cal = 16'b0000010000011100;
            15'd10916: log10_cal = 16'b0000010000011100;
            15'd10917: log10_cal = 16'b0000010000011100;
            15'd10918: log10_cal = 16'b0000010000011100;
            15'd10919: log10_cal = 16'b0000010000011100;
            15'd10920: log10_cal = 16'b0000010000011100;
            15'd10921: log10_cal = 16'b0000010000011100;
            15'd10922: log10_cal = 16'b0000010000011100;
            15'd10923: log10_cal = 16'b0000010000011100;
            15'd10924: log10_cal = 16'b0000010000011100;
            15'd10925: log10_cal = 16'b0000010000011100;
            15'd10926: log10_cal = 16'b0000010000011100;
            15'd10927: log10_cal = 16'b0000010000011100;
            15'd10928: log10_cal = 16'b0000010000011100;
            15'd10929: log10_cal = 16'b0000010000011100;
            15'd10930: log10_cal = 16'b0000010000011100;
            15'd10931: log10_cal = 16'b0000010000011101;
            15'd10932: log10_cal = 16'b0000010000011101;
            15'd10933: log10_cal = 16'b0000010000011101;
            15'd10934: log10_cal = 16'b0000010000011101;
            15'd10935: log10_cal = 16'b0000010000011101;
            15'd10936: log10_cal = 16'b0000010000011101;
            15'd10937: log10_cal = 16'b0000010000011101;
            15'd10938: log10_cal = 16'b0000010000011101;
            15'd10939: log10_cal = 16'b0000010000011101;
            15'd10940: log10_cal = 16'b0000010000011101;
            15'd10941: log10_cal = 16'b0000010000011101;
            15'd10942: log10_cal = 16'b0000010000011101;
            15'd10943: log10_cal = 16'b0000010000011101;
            15'd10944: log10_cal = 16'b0000010000011101;
            15'd10945: log10_cal = 16'b0000010000011101;
            15'd10946: log10_cal = 16'b0000010000011101;
            15'd10947: log10_cal = 16'b0000010000011101;
            15'd10948: log10_cal = 16'b0000010000011101;
            15'd10949: log10_cal = 16'b0000010000011101;
            15'd10950: log10_cal = 16'b0000010000011101;
            15'd10951: log10_cal = 16'b0000010000011101;
            15'd10952: log10_cal = 16'b0000010000011101;
            15'd10953: log10_cal = 16'b0000010000011101;
            15'd10954: log10_cal = 16'b0000010000011101;
            15'd10955: log10_cal = 16'b0000010000011110;
            15'd10956: log10_cal = 16'b0000010000011110;
            15'd10957: log10_cal = 16'b0000010000011110;
            15'd10958: log10_cal = 16'b0000010000011110;
            15'd10959: log10_cal = 16'b0000010000011110;
            15'd10960: log10_cal = 16'b0000010000011110;
            15'd10961: log10_cal = 16'b0000010000011110;
            15'd10962: log10_cal = 16'b0000010000011110;
            15'd10963: log10_cal = 16'b0000010000011110;
            15'd10964: log10_cal = 16'b0000010000011110;
            15'd10965: log10_cal = 16'b0000010000011110;
            15'd10966: log10_cal = 16'b0000010000011110;
            15'd10967: log10_cal = 16'b0000010000011110;
            15'd10968: log10_cal = 16'b0000010000011110;
            15'd10969: log10_cal = 16'b0000010000011110;
            15'd10970: log10_cal = 16'b0000010000011110;
            15'd10971: log10_cal = 16'b0000010000011110;
            15'd10972: log10_cal = 16'b0000010000011110;
            15'd10973: log10_cal = 16'b0000010000011110;
            15'd10974: log10_cal = 16'b0000010000011110;
            15'd10975: log10_cal = 16'b0000010000011110;
            15'd10976: log10_cal = 16'b0000010000011110;
            15'd10977: log10_cal = 16'b0000010000011110;
            15'd10978: log10_cal = 16'b0000010000011110;
            15'd10979: log10_cal = 16'b0000010000011110;
            15'd10980: log10_cal = 16'b0000010000011111;
            15'd10981: log10_cal = 16'b0000010000011111;
            15'd10982: log10_cal = 16'b0000010000011111;
            15'd10983: log10_cal = 16'b0000010000011111;
            15'd10984: log10_cal = 16'b0000010000011111;
            15'd10985: log10_cal = 16'b0000010000011111;
            15'd10986: log10_cal = 16'b0000010000011111;
            15'd10987: log10_cal = 16'b0000010000011111;
            15'd10988: log10_cal = 16'b0000010000011111;
            15'd10989: log10_cal = 16'b0000010000011111;
            15'd10990: log10_cal = 16'b0000010000011111;
            15'd10991: log10_cal = 16'b0000010000011111;
            15'd10992: log10_cal = 16'b0000010000011111;
            15'd10993: log10_cal = 16'b0000010000011111;
            15'd10994: log10_cal = 16'b0000010000011111;
            15'd10995: log10_cal = 16'b0000010000011111;
            15'd10996: log10_cal = 16'b0000010000011111;
            15'd10997: log10_cal = 16'b0000010000011111;
            15'd10998: log10_cal = 16'b0000010000011111;
            15'd10999: log10_cal = 16'b0000010000011111;
            15'd11000: log10_cal = 16'b0000010000011111;
            15'd11001: log10_cal = 16'b0000010000011111;
            15'd11002: log10_cal = 16'b0000010000011111;
            15'd11003: log10_cal = 16'b0000010000011111;
            15'd11004: log10_cal = 16'b0000010000100000;
            15'd11005: log10_cal = 16'b0000010000100000;
            15'd11006: log10_cal = 16'b0000010000100000;
            15'd11007: log10_cal = 16'b0000010000100000;
            15'd11008: log10_cal = 16'b0000010000100000;
            15'd11009: log10_cal = 16'b0000010000100000;
            15'd11010: log10_cal = 16'b0000010000100000;
            15'd11011: log10_cal = 16'b0000010000100000;
            15'd11012: log10_cal = 16'b0000010000100000;
            15'd11013: log10_cal = 16'b0000010000100000;
            15'd11014: log10_cal = 16'b0000010000100000;
            15'd11015: log10_cal = 16'b0000010000100000;
            15'd11016: log10_cal = 16'b0000010000100000;
            15'd11017: log10_cal = 16'b0000010000100000;
            15'd11018: log10_cal = 16'b0000010000100000;
            15'd11019: log10_cal = 16'b0000010000100000;
            15'd11020: log10_cal = 16'b0000010000100000;
            15'd11021: log10_cal = 16'b0000010000100000;
            15'd11022: log10_cal = 16'b0000010000100000;
            15'd11023: log10_cal = 16'b0000010000100000;
            15'd11024: log10_cal = 16'b0000010000100000;
            15'd11025: log10_cal = 16'b0000010000100000;
            15'd11026: log10_cal = 16'b0000010000100000;
            15'd11027: log10_cal = 16'b0000010000100000;
            15'd11028: log10_cal = 16'b0000010000100000;
            15'd11029: log10_cal = 16'b0000010000100001;
            15'd11030: log10_cal = 16'b0000010000100001;
            15'd11031: log10_cal = 16'b0000010000100001;
            15'd11032: log10_cal = 16'b0000010000100001;
            15'd11033: log10_cal = 16'b0000010000100001;
            15'd11034: log10_cal = 16'b0000010000100001;
            15'd11035: log10_cal = 16'b0000010000100001;
            15'd11036: log10_cal = 16'b0000010000100001;
            15'd11037: log10_cal = 16'b0000010000100001;
            15'd11038: log10_cal = 16'b0000010000100001;
            15'd11039: log10_cal = 16'b0000010000100001;
            15'd11040: log10_cal = 16'b0000010000100001;
            15'd11041: log10_cal = 16'b0000010000100001;
            15'd11042: log10_cal = 16'b0000010000100001;
            15'd11043: log10_cal = 16'b0000010000100001;
            15'd11044: log10_cal = 16'b0000010000100001;
            15'd11045: log10_cal = 16'b0000010000100001;
            15'd11046: log10_cal = 16'b0000010000100001;
            15'd11047: log10_cal = 16'b0000010000100001;
            15'd11048: log10_cal = 16'b0000010000100001;
            15'd11049: log10_cal = 16'b0000010000100001;
            15'd11050: log10_cal = 16'b0000010000100001;
            15'd11051: log10_cal = 16'b0000010000100001;
            15'd11052: log10_cal = 16'b0000010000100001;
            15'd11053: log10_cal = 16'b0000010000100001;
            15'd11054: log10_cal = 16'b0000010000100010;
            15'd11055: log10_cal = 16'b0000010000100010;
            15'd11056: log10_cal = 16'b0000010000100010;
            15'd11057: log10_cal = 16'b0000010000100010;
            15'd11058: log10_cal = 16'b0000010000100010;
            15'd11059: log10_cal = 16'b0000010000100010;
            15'd11060: log10_cal = 16'b0000010000100010;
            15'd11061: log10_cal = 16'b0000010000100010;
            15'd11062: log10_cal = 16'b0000010000100010;
            15'd11063: log10_cal = 16'b0000010000100010;
            15'd11064: log10_cal = 16'b0000010000100010;
            15'd11065: log10_cal = 16'b0000010000100010;
            15'd11066: log10_cal = 16'b0000010000100010;
            15'd11067: log10_cal = 16'b0000010000100010;
            15'd11068: log10_cal = 16'b0000010000100010;
            15'd11069: log10_cal = 16'b0000010000100010;
            15'd11070: log10_cal = 16'b0000010000100010;
            15'd11071: log10_cal = 16'b0000010000100010;
            15'd11072: log10_cal = 16'b0000010000100010;
            15'd11073: log10_cal = 16'b0000010000100010;
            15'd11074: log10_cal = 16'b0000010000100010;
            15'd11075: log10_cal = 16'b0000010000100010;
            15'd11076: log10_cal = 16'b0000010000100010;
            15'd11077: log10_cal = 16'b0000010000100010;
            15'd11078: log10_cal = 16'b0000010000100010;
            15'd11079: log10_cal = 16'b0000010000100011;
            15'd11080: log10_cal = 16'b0000010000100011;
            15'd11081: log10_cal = 16'b0000010000100011;
            15'd11082: log10_cal = 16'b0000010000100011;
            15'd11083: log10_cal = 16'b0000010000100011;
            15'd11084: log10_cal = 16'b0000010000100011;
            15'd11085: log10_cal = 16'b0000010000100011;
            15'd11086: log10_cal = 16'b0000010000100011;
            15'd11087: log10_cal = 16'b0000010000100011;
            15'd11088: log10_cal = 16'b0000010000100011;
            15'd11089: log10_cal = 16'b0000010000100011;
            15'd11090: log10_cal = 16'b0000010000100011;
            15'd11091: log10_cal = 16'b0000010000100011;
            15'd11092: log10_cal = 16'b0000010000100011;
            15'd11093: log10_cal = 16'b0000010000100011;
            15'd11094: log10_cal = 16'b0000010000100011;
            15'd11095: log10_cal = 16'b0000010000100011;
            15'd11096: log10_cal = 16'b0000010000100011;
            15'd11097: log10_cal = 16'b0000010000100011;
            15'd11098: log10_cal = 16'b0000010000100011;
            15'd11099: log10_cal = 16'b0000010000100011;
            15'd11100: log10_cal = 16'b0000010000100011;
            15'd11101: log10_cal = 16'b0000010000100011;
            15'd11102: log10_cal = 16'b0000010000100011;
            15'd11103: log10_cal = 16'b0000010000100011;
            15'd11104: log10_cal = 16'b0000010000100100;
            15'd11105: log10_cal = 16'b0000010000100100;
            15'd11106: log10_cal = 16'b0000010000100100;
            15'd11107: log10_cal = 16'b0000010000100100;
            15'd11108: log10_cal = 16'b0000010000100100;
            15'd11109: log10_cal = 16'b0000010000100100;
            15'd11110: log10_cal = 16'b0000010000100100;
            15'd11111: log10_cal = 16'b0000010000100100;
            15'd11112: log10_cal = 16'b0000010000100100;
            15'd11113: log10_cal = 16'b0000010000100100;
            15'd11114: log10_cal = 16'b0000010000100100;
            15'd11115: log10_cal = 16'b0000010000100100;
            15'd11116: log10_cal = 16'b0000010000100100;
            15'd11117: log10_cal = 16'b0000010000100100;
            15'd11118: log10_cal = 16'b0000010000100100;
            15'd11119: log10_cal = 16'b0000010000100100;
            15'd11120: log10_cal = 16'b0000010000100100;
            15'd11121: log10_cal = 16'b0000010000100100;
            15'd11122: log10_cal = 16'b0000010000100100;
            15'd11123: log10_cal = 16'b0000010000100100;
            15'd11124: log10_cal = 16'b0000010000100100;
            15'd11125: log10_cal = 16'b0000010000100100;
            15'd11126: log10_cal = 16'b0000010000100100;
            15'd11127: log10_cal = 16'b0000010000100100;
            15'd11128: log10_cal = 16'b0000010000100100;
            15'd11129: log10_cal = 16'b0000010000100101;
            15'd11130: log10_cal = 16'b0000010000100101;
            15'd11131: log10_cal = 16'b0000010000100101;
            15'd11132: log10_cal = 16'b0000010000100101;
            15'd11133: log10_cal = 16'b0000010000100101;
            15'd11134: log10_cal = 16'b0000010000100101;
            15'd11135: log10_cal = 16'b0000010000100101;
            15'd11136: log10_cal = 16'b0000010000100101;
            15'd11137: log10_cal = 16'b0000010000100101;
            15'd11138: log10_cal = 16'b0000010000100101;
            15'd11139: log10_cal = 16'b0000010000100101;
            15'd11140: log10_cal = 16'b0000010000100101;
            15'd11141: log10_cal = 16'b0000010000100101;
            15'd11142: log10_cal = 16'b0000010000100101;
            15'd11143: log10_cal = 16'b0000010000100101;
            15'd11144: log10_cal = 16'b0000010000100101;
            15'd11145: log10_cal = 16'b0000010000100101;
            15'd11146: log10_cal = 16'b0000010000100101;
            15'd11147: log10_cal = 16'b0000010000100101;
            15'd11148: log10_cal = 16'b0000010000100101;
            15'd11149: log10_cal = 16'b0000010000100101;
            15'd11150: log10_cal = 16'b0000010000100101;
            15'd11151: log10_cal = 16'b0000010000100101;
            15'd11152: log10_cal = 16'b0000010000100101;
            15'd11153: log10_cal = 16'b0000010000100101;
            15'd11154: log10_cal = 16'b0000010000100110;
            15'd11155: log10_cal = 16'b0000010000100110;
            15'd11156: log10_cal = 16'b0000010000100110;
            15'd11157: log10_cal = 16'b0000010000100110;
            15'd11158: log10_cal = 16'b0000010000100110;
            15'd11159: log10_cal = 16'b0000010000100110;
            15'd11160: log10_cal = 16'b0000010000100110;
            15'd11161: log10_cal = 16'b0000010000100110;
            15'd11162: log10_cal = 16'b0000010000100110;
            15'd11163: log10_cal = 16'b0000010000100110;
            15'd11164: log10_cal = 16'b0000010000100110;
            15'd11165: log10_cal = 16'b0000010000100110;
            15'd11166: log10_cal = 16'b0000010000100110;
            15'd11167: log10_cal = 16'b0000010000100110;
            15'd11168: log10_cal = 16'b0000010000100110;
            15'd11169: log10_cal = 16'b0000010000100110;
            15'd11170: log10_cal = 16'b0000010000100110;
            15'd11171: log10_cal = 16'b0000010000100110;
            15'd11172: log10_cal = 16'b0000010000100110;
            15'd11173: log10_cal = 16'b0000010000100110;
            15'd11174: log10_cal = 16'b0000010000100110;
            15'd11175: log10_cal = 16'b0000010000100110;
            15'd11176: log10_cal = 16'b0000010000100110;
            15'd11177: log10_cal = 16'b0000010000100110;
            15'd11178: log10_cal = 16'b0000010000100110;
            15'd11179: log10_cal = 16'b0000010000100111;
            15'd11180: log10_cal = 16'b0000010000100111;
            15'd11181: log10_cal = 16'b0000010000100111;
            15'd11182: log10_cal = 16'b0000010000100111;
            15'd11183: log10_cal = 16'b0000010000100111;
            15'd11184: log10_cal = 16'b0000010000100111;
            15'd11185: log10_cal = 16'b0000010000100111;
            15'd11186: log10_cal = 16'b0000010000100111;
            15'd11187: log10_cal = 16'b0000010000100111;
            15'd11188: log10_cal = 16'b0000010000100111;
            15'd11189: log10_cal = 16'b0000010000100111;
            15'd11190: log10_cal = 16'b0000010000100111;
            15'd11191: log10_cal = 16'b0000010000100111;
            15'd11192: log10_cal = 16'b0000010000100111;
            15'd11193: log10_cal = 16'b0000010000100111;
            15'd11194: log10_cal = 16'b0000010000100111;
            15'd11195: log10_cal = 16'b0000010000100111;
            15'd11196: log10_cal = 16'b0000010000100111;
            15'd11197: log10_cal = 16'b0000010000100111;
            15'd11198: log10_cal = 16'b0000010000100111;
            15'd11199: log10_cal = 16'b0000010000100111;
            15'd11200: log10_cal = 16'b0000010000100111;
            15'd11201: log10_cal = 16'b0000010000100111;
            15'd11202: log10_cal = 16'b0000010000100111;
            15'd11203: log10_cal = 16'b0000010000100111;
            15'd11204: log10_cal = 16'b0000010000101000;
            15'd11205: log10_cal = 16'b0000010000101000;
            15'd11206: log10_cal = 16'b0000010000101000;
            15'd11207: log10_cal = 16'b0000010000101000;
            15'd11208: log10_cal = 16'b0000010000101000;
            15'd11209: log10_cal = 16'b0000010000101000;
            15'd11210: log10_cal = 16'b0000010000101000;
            15'd11211: log10_cal = 16'b0000010000101000;
            15'd11212: log10_cal = 16'b0000010000101000;
            15'd11213: log10_cal = 16'b0000010000101000;
            15'd11214: log10_cal = 16'b0000010000101000;
            15'd11215: log10_cal = 16'b0000010000101000;
            15'd11216: log10_cal = 16'b0000010000101000;
            15'd11217: log10_cal = 16'b0000010000101000;
            15'd11218: log10_cal = 16'b0000010000101000;
            15'd11219: log10_cal = 16'b0000010000101000;
            15'd11220: log10_cal = 16'b0000010000101000;
            15'd11221: log10_cal = 16'b0000010000101000;
            15'd11222: log10_cal = 16'b0000010000101000;
            15'd11223: log10_cal = 16'b0000010000101000;
            15'd11224: log10_cal = 16'b0000010000101000;
            15'd11225: log10_cal = 16'b0000010000101000;
            15'd11226: log10_cal = 16'b0000010000101000;
            15'd11227: log10_cal = 16'b0000010000101000;
            15'd11228: log10_cal = 16'b0000010000101000;
            15'd11229: log10_cal = 16'b0000010000101001;
            15'd11230: log10_cal = 16'b0000010000101001;
            15'd11231: log10_cal = 16'b0000010000101001;
            15'd11232: log10_cal = 16'b0000010000101001;
            15'd11233: log10_cal = 16'b0000010000101001;
            15'd11234: log10_cal = 16'b0000010000101001;
            15'd11235: log10_cal = 16'b0000010000101001;
            15'd11236: log10_cal = 16'b0000010000101001;
            15'd11237: log10_cal = 16'b0000010000101001;
            15'd11238: log10_cal = 16'b0000010000101001;
            15'd11239: log10_cal = 16'b0000010000101001;
            15'd11240: log10_cal = 16'b0000010000101001;
            15'd11241: log10_cal = 16'b0000010000101001;
            15'd11242: log10_cal = 16'b0000010000101001;
            15'd11243: log10_cal = 16'b0000010000101001;
            15'd11244: log10_cal = 16'b0000010000101001;
            15'd11245: log10_cal = 16'b0000010000101001;
            15'd11246: log10_cal = 16'b0000010000101001;
            15'd11247: log10_cal = 16'b0000010000101001;
            15'd11248: log10_cal = 16'b0000010000101001;
            15'd11249: log10_cal = 16'b0000010000101001;
            15'd11250: log10_cal = 16'b0000010000101001;
            15'd11251: log10_cal = 16'b0000010000101001;
            15'd11252: log10_cal = 16'b0000010000101001;
            15'd11253: log10_cal = 16'b0000010000101001;
            15'd11254: log10_cal = 16'b0000010000101001;
            15'd11255: log10_cal = 16'b0000010000101010;
            15'd11256: log10_cal = 16'b0000010000101010;
            15'd11257: log10_cal = 16'b0000010000101010;
            15'd11258: log10_cal = 16'b0000010000101010;
            15'd11259: log10_cal = 16'b0000010000101010;
            15'd11260: log10_cal = 16'b0000010000101010;
            15'd11261: log10_cal = 16'b0000010000101010;
            15'd11262: log10_cal = 16'b0000010000101010;
            15'd11263: log10_cal = 16'b0000010000101010;
            15'd11264: log10_cal = 16'b0000010000101010;
            15'd11265: log10_cal = 16'b0000010000101010;
            15'd11266: log10_cal = 16'b0000010000101010;
            15'd11267: log10_cal = 16'b0000010000101010;
            15'd11268: log10_cal = 16'b0000010000101010;
            15'd11269: log10_cal = 16'b0000010000101010;
            15'd11270: log10_cal = 16'b0000010000101010;
            15'd11271: log10_cal = 16'b0000010000101010;
            15'd11272: log10_cal = 16'b0000010000101010;
            15'd11273: log10_cal = 16'b0000010000101010;
            15'd11274: log10_cal = 16'b0000010000101010;
            15'd11275: log10_cal = 16'b0000010000101010;
            15'd11276: log10_cal = 16'b0000010000101010;
            15'd11277: log10_cal = 16'b0000010000101010;
            15'd11278: log10_cal = 16'b0000010000101010;
            15'd11279: log10_cal = 16'b0000010000101010;
            15'd11280: log10_cal = 16'b0000010000101011;
            15'd11281: log10_cal = 16'b0000010000101011;
            15'd11282: log10_cal = 16'b0000010000101011;
            15'd11283: log10_cal = 16'b0000010000101011;
            15'd11284: log10_cal = 16'b0000010000101011;
            15'd11285: log10_cal = 16'b0000010000101011;
            15'd11286: log10_cal = 16'b0000010000101011;
            15'd11287: log10_cal = 16'b0000010000101011;
            15'd11288: log10_cal = 16'b0000010000101011;
            15'd11289: log10_cal = 16'b0000010000101011;
            15'd11290: log10_cal = 16'b0000010000101011;
            15'd11291: log10_cal = 16'b0000010000101011;
            15'd11292: log10_cal = 16'b0000010000101011;
            15'd11293: log10_cal = 16'b0000010000101011;
            15'd11294: log10_cal = 16'b0000010000101011;
            15'd11295: log10_cal = 16'b0000010000101011;
            15'd11296: log10_cal = 16'b0000010000101011;
            15'd11297: log10_cal = 16'b0000010000101011;
            15'd11298: log10_cal = 16'b0000010000101011;
            15'd11299: log10_cal = 16'b0000010000101011;
            15'd11300: log10_cal = 16'b0000010000101011;
            15'd11301: log10_cal = 16'b0000010000101011;
            15'd11302: log10_cal = 16'b0000010000101011;
            15'd11303: log10_cal = 16'b0000010000101011;
            15'd11304: log10_cal = 16'b0000010000101011;
            15'd11305: log10_cal = 16'b0000010000101100;
            15'd11306: log10_cal = 16'b0000010000101100;
            15'd11307: log10_cal = 16'b0000010000101100;
            15'd11308: log10_cal = 16'b0000010000101100;
            15'd11309: log10_cal = 16'b0000010000101100;
            15'd11310: log10_cal = 16'b0000010000101100;
            15'd11311: log10_cal = 16'b0000010000101100;
            15'd11312: log10_cal = 16'b0000010000101100;
            15'd11313: log10_cal = 16'b0000010000101100;
            15'd11314: log10_cal = 16'b0000010000101100;
            15'd11315: log10_cal = 16'b0000010000101100;
            15'd11316: log10_cal = 16'b0000010000101100;
            15'd11317: log10_cal = 16'b0000010000101100;
            15'd11318: log10_cal = 16'b0000010000101100;
            15'd11319: log10_cal = 16'b0000010000101100;
            15'd11320: log10_cal = 16'b0000010000101100;
            15'd11321: log10_cal = 16'b0000010000101100;
            15'd11322: log10_cal = 16'b0000010000101100;
            15'd11323: log10_cal = 16'b0000010000101100;
            15'd11324: log10_cal = 16'b0000010000101100;
            15'd11325: log10_cal = 16'b0000010000101100;
            15'd11326: log10_cal = 16'b0000010000101100;
            15'd11327: log10_cal = 16'b0000010000101100;
            15'd11328: log10_cal = 16'b0000010000101100;
            15'd11329: log10_cal = 16'b0000010000101100;
            15'd11330: log10_cal = 16'b0000010000101100;
            15'd11331: log10_cal = 16'b0000010000101101;
            15'd11332: log10_cal = 16'b0000010000101101;
            15'd11333: log10_cal = 16'b0000010000101101;
            15'd11334: log10_cal = 16'b0000010000101101;
            15'd11335: log10_cal = 16'b0000010000101101;
            15'd11336: log10_cal = 16'b0000010000101101;
            15'd11337: log10_cal = 16'b0000010000101101;
            15'd11338: log10_cal = 16'b0000010000101101;
            15'd11339: log10_cal = 16'b0000010000101101;
            15'd11340: log10_cal = 16'b0000010000101101;
            15'd11341: log10_cal = 16'b0000010000101101;
            15'd11342: log10_cal = 16'b0000010000101101;
            15'd11343: log10_cal = 16'b0000010000101101;
            15'd11344: log10_cal = 16'b0000010000101101;
            15'd11345: log10_cal = 16'b0000010000101101;
            15'd11346: log10_cal = 16'b0000010000101101;
            15'd11347: log10_cal = 16'b0000010000101101;
            15'd11348: log10_cal = 16'b0000010000101101;
            15'd11349: log10_cal = 16'b0000010000101101;
            15'd11350: log10_cal = 16'b0000010000101101;
            15'd11351: log10_cal = 16'b0000010000101101;
            15'd11352: log10_cal = 16'b0000010000101101;
            15'd11353: log10_cal = 16'b0000010000101101;
            15'd11354: log10_cal = 16'b0000010000101101;
            15'd11355: log10_cal = 16'b0000010000101101;
            15'd11356: log10_cal = 16'b0000010000101110;
            15'd11357: log10_cal = 16'b0000010000101110;
            15'd11358: log10_cal = 16'b0000010000101110;
            15'd11359: log10_cal = 16'b0000010000101110;
            15'd11360: log10_cal = 16'b0000010000101110;
            15'd11361: log10_cal = 16'b0000010000101110;
            15'd11362: log10_cal = 16'b0000010000101110;
            15'd11363: log10_cal = 16'b0000010000101110;
            15'd11364: log10_cal = 16'b0000010000101110;
            15'd11365: log10_cal = 16'b0000010000101110;
            15'd11366: log10_cal = 16'b0000010000101110;
            15'd11367: log10_cal = 16'b0000010000101110;
            15'd11368: log10_cal = 16'b0000010000101110;
            15'd11369: log10_cal = 16'b0000010000101110;
            15'd11370: log10_cal = 16'b0000010000101110;
            15'd11371: log10_cal = 16'b0000010000101110;
            15'd11372: log10_cal = 16'b0000010000101110;
            15'd11373: log10_cal = 16'b0000010000101110;
            15'd11374: log10_cal = 16'b0000010000101110;
            15'd11375: log10_cal = 16'b0000010000101110;
            15'd11376: log10_cal = 16'b0000010000101110;
            15'd11377: log10_cal = 16'b0000010000101110;
            15'd11378: log10_cal = 16'b0000010000101110;
            15'd11379: log10_cal = 16'b0000010000101110;
            15'd11380: log10_cal = 16'b0000010000101110;
            15'd11381: log10_cal = 16'b0000010000101110;
            15'd11382: log10_cal = 16'b0000010000101111;
            15'd11383: log10_cal = 16'b0000010000101111;
            15'd11384: log10_cal = 16'b0000010000101111;
            15'd11385: log10_cal = 16'b0000010000101111;
            15'd11386: log10_cal = 16'b0000010000101111;
            15'd11387: log10_cal = 16'b0000010000101111;
            15'd11388: log10_cal = 16'b0000010000101111;
            15'd11389: log10_cal = 16'b0000010000101111;
            15'd11390: log10_cal = 16'b0000010000101111;
            15'd11391: log10_cal = 16'b0000010000101111;
            15'd11392: log10_cal = 16'b0000010000101111;
            15'd11393: log10_cal = 16'b0000010000101111;
            15'd11394: log10_cal = 16'b0000010000101111;
            15'd11395: log10_cal = 16'b0000010000101111;
            15'd11396: log10_cal = 16'b0000010000101111;
            15'd11397: log10_cal = 16'b0000010000101111;
            15'd11398: log10_cal = 16'b0000010000101111;
            15'd11399: log10_cal = 16'b0000010000101111;
            15'd11400: log10_cal = 16'b0000010000101111;
            15'd11401: log10_cal = 16'b0000010000101111;
            15'd11402: log10_cal = 16'b0000010000101111;
            15'd11403: log10_cal = 16'b0000010000101111;
            15'd11404: log10_cal = 16'b0000010000101111;
            15'd11405: log10_cal = 16'b0000010000101111;
            15'd11406: log10_cal = 16'b0000010000101111;
            15'd11407: log10_cal = 16'b0000010000101111;
            15'd11408: log10_cal = 16'b0000010000110000;
            15'd11409: log10_cal = 16'b0000010000110000;
            15'd11410: log10_cal = 16'b0000010000110000;
            15'd11411: log10_cal = 16'b0000010000110000;
            15'd11412: log10_cal = 16'b0000010000110000;
            15'd11413: log10_cal = 16'b0000010000110000;
            15'd11414: log10_cal = 16'b0000010000110000;
            15'd11415: log10_cal = 16'b0000010000110000;
            15'd11416: log10_cal = 16'b0000010000110000;
            15'd11417: log10_cal = 16'b0000010000110000;
            15'd11418: log10_cal = 16'b0000010000110000;
            15'd11419: log10_cal = 16'b0000010000110000;
            15'd11420: log10_cal = 16'b0000010000110000;
            15'd11421: log10_cal = 16'b0000010000110000;
            15'd11422: log10_cal = 16'b0000010000110000;
            15'd11423: log10_cal = 16'b0000010000110000;
            15'd11424: log10_cal = 16'b0000010000110000;
            15'd11425: log10_cal = 16'b0000010000110000;
            15'd11426: log10_cal = 16'b0000010000110000;
            15'd11427: log10_cal = 16'b0000010000110000;
            15'd11428: log10_cal = 16'b0000010000110000;
            15'd11429: log10_cal = 16'b0000010000110000;
            15'd11430: log10_cal = 16'b0000010000110000;
            15'd11431: log10_cal = 16'b0000010000110000;
            15'd11432: log10_cal = 16'b0000010000110000;
            15'd11433: log10_cal = 16'b0000010000110001;
            15'd11434: log10_cal = 16'b0000010000110001;
            15'd11435: log10_cal = 16'b0000010000110001;
            15'd11436: log10_cal = 16'b0000010000110001;
            15'd11437: log10_cal = 16'b0000010000110001;
            15'd11438: log10_cal = 16'b0000010000110001;
            15'd11439: log10_cal = 16'b0000010000110001;
            15'd11440: log10_cal = 16'b0000010000110001;
            15'd11441: log10_cal = 16'b0000010000110001;
            15'd11442: log10_cal = 16'b0000010000110001;
            15'd11443: log10_cal = 16'b0000010000110001;
            15'd11444: log10_cal = 16'b0000010000110001;
            15'd11445: log10_cal = 16'b0000010000110001;
            15'd11446: log10_cal = 16'b0000010000110001;
            15'd11447: log10_cal = 16'b0000010000110001;
            15'd11448: log10_cal = 16'b0000010000110001;
            15'd11449: log10_cal = 16'b0000010000110001;
            15'd11450: log10_cal = 16'b0000010000110001;
            15'd11451: log10_cal = 16'b0000010000110001;
            15'd11452: log10_cal = 16'b0000010000110001;
            15'd11453: log10_cal = 16'b0000010000110001;
            15'd11454: log10_cal = 16'b0000010000110001;
            15'd11455: log10_cal = 16'b0000010000110001;
            15'd11456: log10_cal = 16'b0000010000110001;
            15'd11457: log10_cal = 16'b0000010000110001;
            15'd11458: log10_cal = 16'b0000010000110001;
            15'd11459: log10_cal = 16'b0000010000110010;
            15'd11460: log10_cal = 16'b0000010000110010;
            15'd11461: log10_cal = 16'b0000010000110010;
            15'd11462: log10_cal = 16'b0000010000110010;
            15'd11463: log10_cal = 16'b0000010000110010;
            15'd11464: log10_cal = 16'b0000010000110010;
            15'd11465: log10_cal = 16'b0000010000110010;
            15'd11466: log10_cal = 16'b0000010000110010;
            15'd11467: log10_cal = 16'b0000010000110010;
            15'd11468: log10_cal = 16'b0000010000110010;
            15'd11469: log10_cal = 16'b0000010000110010;
            15'd11470: log10_cal = 16'b0000010000110010;
            15'd11471: log10_cal = 16'b0000010000110010;
            15'd11472: log10_cal = 16'b0000010000110010;
            15'd11473: log10_cal = 16'b0000010000110010;
            15'd11474: log10_cal = 16'b0000010000110010;
            15'd11475: log10_cal = 16'b0000010000110010;
            15'd11476: log10_cal = 16'b0000010000110010;
            15'd11477: log10_cal = 16'b0000010000110010;
            15'd11478: log10_cal = 16'b0000010000110010;
            15'd11479: log10_cal = 16'b0000010000110010;
            15'd11480: log10_cal = 16'b0000010000110010;
            15'd11481: log10_cal = 16'b0000010000110010;
            15'd11482: log10_cal = 16'b0000010000110010;
            15'd11483: log10_cal = 16'b0000010000110010;
            15'd11484: log10_cal = 16'b0000010000110010;
            15'd11485: log10_cal = 16'b0000010000110011;
            15'd11486: log10_cal = 16'b0000010000110011;
            15'd11487: log10_cal = 16'b0000010000110011;
            15'd11488: log10_cal = 16'b0000010000110011;
            15'd11489: log10_cal = 16'b0000010000110011;
            15'd11490: log10_cal = 16'b0000010000110011;
            15'd11491: log10_cal = 16'b0000010000110011;
            15'd11492: log10_cal = 16'b0000010000110011;
            15'd11493: log10_cal = 16'b0000010000110011;
            15'd11494: log10_cal = 16'b0000010000110011;
            15'd11495: log10_cal = 16'b0000010000110011;
            15'd11496: log10_cal = 16'b0000010000110011;
            15'd11497: log10_cal = 16'b0000010000110011;
            15'd11498: log10_cal = 16'b0000010000110011;
            15'd11499: log10_cal = 16'b0000010000110011;
            15'd11500: log10_cal = 16'b0000010000110011;
            15'd11501: log10_cal = 16'b0000010000110011;
            15'd11502: log10_cal = 16'b0000010000110011;
            15'd11503: log10_cal = 16'b0000010000110011;
            15'd11504: log10_cal = 16'b0000010000110011;
            15'd11505: log10_cal = 16'b0000010000110011;
            15'd11506: log10_cal = 16'b0000010000110011;
            15'd11507: log10_cal = 16'b0000010000110011;
            15'd11508: log10_cal = 16'b0000010000110011;
            15'd11509: log10_cal = 16'b0000010000110011;
            15'd11510: log10_cal = 16'b0000010000110011;
            15'd11511: log10_cal = 16'b0000010000110100;
            15'd11512: log10_cal = 16'b0000010000110100;
            15'd11513: log10_cal = 16'b0000010000110100;
            15'd11514: log10_cal = 16'b0000010000110100;
            15'd11515: log10_cal = 16'b0000010000110100;
            15'd11516: log10_cal = 16'b0000010000110100;
            15'd11517: log10_cal = 16'b0000010000110100;
            15'd11518: log10_cal = 16'b0000010000110100;
            15'd11519: log10_cal = 16'b0000010000110100;
            15'd11520: log10_cal = 16'b0000010000110100;
            15'd11521: log10_cal = 16'b0000010000110100;
            15'd11522: log10_cal = 16'b0000010000110100;
            15'd11523: log10_cal = 16'b0000010000110100;
            15'd11524: log10_cal = 16'b0000010000110100;
            15'd11525: log10_cal = 16'b0000010000110100;
            15'd11526: log10_cal = 16'b0000010000110100;
            15'd11527: log10_cal = 16'b0000010000110100;
            15'd11528: log10_cal = 16'b0000010000110100;
            15'd11529: log10_cal = 16'b0000010000110100;
            15'd11530: log10_cal = 16'b0000010000110100;
            15'd11531: log10_cal = 16'b0000010000110100;
            15'd11532: log10_cal = 16'b0000010000110100;
            15'd11533: log10_cal = 16'b0000010000110100;
            15'd11534: log10_cal = 16'b0000010000110100;
            15'd11535: log10_cal = 16'b0000010000110100;
            15'd11536: log10_cal = 16'b0000010000110100;
            15'd11537: log10_cal = 16'b0000010000110101;
            15'd11538: log10_cal = 16'b0000010000110101;
            15'd11539: log10_cal = 16'b0000010000110101;
            15'd11540: log10_cal = 16'b0000010000110101;
            15'd11541: log10_cal = 16'b0000010000110101;
            15'd11542: log10_cal = 16'b0000010000110101;
            15'd11543: log10_cal = 16'b0000010000110101;
            15'd11544: log10_cal = 16'b0000010000110101;
            15'd11545: log10_cal = 16'b0000010000110101;
            15'd11546: log10_cal = 16'b0000010000110101;
            15'd11547: log10_cal = 16'b0000010000110101;
            15'd11548: log10_cal = 16'b0000010000110101;
            15'd11549: log10_cal = 16'b0000010000110101;
            15'd11550: log10_cal = 16'b0000010000110101;
            15'd11551: log10_cal = 16'b0000010000110101;
            15'd11552: log10_cal = 16'b0000010000110101;
            15'd11553: log10_cal = 16'b0000010000110101;
            15'd11554: log10_cal = 16'b0000010000110101;
            15'd11555: log10_cal = 16'b0000010000110101;
            15'd11556: log10_cal = 16'b0000010000110101;
            15'd11557: log10_cal = 16'b0000010000110101;
            15'd11558: log10_cal = 16'b0000010000110101;
            15'd11559: log10_cal = 16'b0000010000110101;
            15'd11560: log10_cal = 16'b0000010000110101;
            15'd11561: log10_cal = 16'b0000010000110101;
            15'd11562: log10_cal = 16'b0000010000110101;
            15'd11563: log10_cal = 16'b0000010000110110;
            15'd11564: log10_cal = 16'b0000010000110110;
            15'd11565: log10_cal = 16'b0000010000110110;
            15'd11566: log10_cal = 16'b0000010000110110;
            15'd11567: log10_cal = 16'b0000010000110110;
            15'd11568: log10_cal = 16'b0000010000110110;
            15'd11569: log10_cal = 16'b0000010000110110;
            15'd11570: log10_cal = 16'b0000010000110110;
            15'd11571: log10_cal = 16'b0000010000110110;
            15'd11572: log10_cal = 16'b0000010000110110;
            15'd11573: log10_cal = 16'b0000010000110110;
            15'd11574: log10_cal = 16'b0000010000110110;
            15'd11575: log10_cal = 16'b0000010000110110;
            15'd11576: log10_cal = 16'b0000010000110110;
            15'd11577: log10_cal = 16'b0000010000110110;
            15'd11578: log10_cal = 16'b0000010000110110;
            15'd11579: log10_cal = 16'b0000010000110110;
            15'd11580: log10_cal = 16'b0000010000110110;
            15'd11581: log10_cal = 16'b0000010000110110;
            15'd11582: log10_cal = 16'b0000010000110110;
            15'd11583: log10_cal = 16'b0000010000110110;
            15'd11584: log10_cal = 16'b0000010000110110;
            15'd11585: log10_cal = 16'b0000010000110110;
            15'd11586: log10_cal = 16'b0000010000110110;
            15'd11587: log10_cal = 16'b0000010000110110;
            15'd11588: log10_cal = 16'b0000010000110110;
            15'd11589: log10_cal = 16'b0000010000110111;
            15'd11590: log10_cal = 16'b0000010000110111;
            15'd11591: log10_cal = 16'b0000010000110111;
            15'd11592: log10_cal = 16'b0000010000110111;
            15'd11593: log10_cal = 16'b0000010000110111;
            15'd11594: log10_cal = 16'b0000010000110111;
            15'd11595: log10_cal = 16'b0000010000110111;
            15'd11596: log10_cal = 16'b0000010000110111;
            15'd11597: log10_cal = 16'b0000010000110111;
            15'd11598: log10_cal = 16'b0000010000110111;
            15'd11599: log10_cal = 16'b0000010000110111;
            15'd11600: log10_cal = 16'b0000010000110111;
            15'd11601: log10_cal = 16'b0000010000110111;
            15'd11602: log10_cal = 16'b0000010000110111;
            15'd11603: log10_cal = 16'b0000010000110111;
            15'd11604: log10_cal = 16'b0000010000110111;
            15'd11605: log10_cal = 16'b0000010000110111;
            15'd11606: log10_cal = 16'b0000010000110111;
            15'd11607: log10_cal = 16'b0000010000110111;
            15'd11608: log10_cal = 16'b0000010000110111;
            15'd11609: log10_cal = 16'b0000010000110111;
            15'd11610: log10_cal = 16'b0000010000110111;
            15'd11611: log10_cal = 16'b0000010000110111;
            15'd11612: log10_cal = 16'b0000010000110111;
            15'd11613: log10_cal = 16'b0000010000110111;
            15'd11614: log10_cal = 16'b0000010000110111;
            15'd11615: log10_cal = 16'b0000010000111000;
            15'd11616: log10_cal = 16'b0000010000111000;
            15'd11617: log10_cal = 16'b0000010000111000;
            15'd11618: log10_cal = 16'b0000010000111000;
            15'd11619: log10_cal = 16'b0000010000111000;
            15'd11620: log10_cal = 16'b0000010000111000;
            15'd11621: log10_cal = 16'b0000010000111000;
            15'd11622: log10_cal = 16'b0000010000111000;
            15'd11623: log10_cal = 16'b0000010000111000;
            15'd11624: log10_cal = 16'b0000010000111000;
            15'd11625: log10_cal = 16'b0000010000111000;
            15'd11626: log10_cal = 16'b0000010000111000;
            15'd11627: log10_cal = 16'b0000010000111000;
            15'd11628: log10_cal = 16'b0000010000111000;
            15'd11629: log10_cal = 16'b0000010000111000;
            15'd11630: log10_cal = 16'b0000010000111000;
            15'd11631: log10_cal = 16'b0000010000111000;
            15'd11632: log10_cal = 16'b0000010000111000;
            15'd11633: log10_cal = 16'b0000010000111000;
            15'd11634: log10_cal = 16'b0000010000111000;
            15'd11635: log10_cal = 16'b0000010000111000;
            15'd11636: log10_cal = 16'b0000010000111000;
            15'd11637: log10_cal = 16'b0000010000111000;
            15'd11638: log10_cal = 16'b0000010000111000;
            15'd11639: log10_cal = 16'b0000010000111000;
            15'd11640: log10_cal = 16'b0000010000111000;
            15'd11641: log10_cal = 16'b0000010000111001;
            15'd11642: log10_cal = 16'b0000010000111001;
            15'd11643: log10_cal = 16'b0000010000111001;
            15'd11644: log10_cal = 16'b0000010000111001;
            15'd11645: log10_cal = 16'b0000010000111001;
            15'd11646: log10_cal = 16'b0000010000111001;
            15'd11647: log10_cal = 16'b0000010000111001;
            15'd11648: log10_cal = 16'b0000010000111001;
            15'd11649: log10_cal = 16'b0000010000111001;
            15'd11650: log10_cal = 16'b0000010000111001;
            15'd11651: log10_cal = 16'b0000010000111001;
            15'd11652: log10_cal = 16'b0000010000111001;
            15'd11653: log10_cal = 16'b0000010000111001;
            15'd11654: log10_cal = 16'b0000010000111001;
            15'd11655: log10_cal = 16'b0000010000111001;
            15'd11656: log10_cal = 16'b0000010000111001;
            15'd11657: log10_cal = 16'b0000010000111001;
            15'd11658: log10_cal = 16'b0000010000111001;
            15'd11659: log10_cal = 16'b0000010000111001;
            15'd11660: log10_cal = 16'b0000010000111001;
            15'd11661: log10_cal = 16'b0000010000111001;
            15'd11662: log10_cal = 16'b0000010000111001;
            15'd11663: log10_cal = 16'b0000010000111001;
            15'd11664: log10_cal = 16'b0000010000111001;
            15'd11665: log10_cal = 16'b0000010000111001;
            15'd11666: log10_cal = 16'b0000010000111001;
            15'd11667: log10_cal = 16'b0000010000111010;
            15'd11668: log10_cal = 16'b0000010000111010;
            15'd11669: log10_cal = 16'b0000010000111010;
            15'd11670: log10_cal = 16'b0000010000111010;
            15'd11671: log10_cal = 16'b0000010000111010;
            15'd11672: log10_cal = 16'b0000010000111010;
            15'd11673: log10_cal = 16'b0000010000111010;
            15'd11674: log10_cal = 16'b0000010000111010;
            15'd11675: log10_cal = 16'b0000010000111010;
            15'd11676: log10_cal = 16'b0000010000111010;
            15'd11677: log10_cal = 16'b0000010000111010;
            15'd11678: log10_cal = 16'b0000010000111010;
            15'd11679: log10_cal = 16'b0000010000111010;
            15'd11680: log10_cal = 16'b0000010000111010;
            15'd11681: log10_cal = 16'b0000010000111010;
            15'd11682: log10_cal = 16'b0000010000111010;
            15'd11683: log10_cal = 16'b0000010000111010;
            15'd11684: log10_cal = 16'b0000010000111010;
            15'd11685: log10_cal = 16'b0000010000111010;
            15'd11686: log10_cal = 16'b0000010000111010;
            15'd11687: log10_cal = 16'b0000010000111010;
            15'd11688: log10_cal = 16'b0000010000111010;
            15'd11689: log10_cal = 16'b0000010000111010;
            15'd11690: log10_cal = 16'b0000010000111010;
            15'd11691: log10_cal = 16'b0000010000111010;
            15'd11692: log10_cal = 16'b0000010000111010;
            15'd11693: log10_cal = 16'b0000010000111011;
            15'd11694: log10_cal = 16'b0000010000111011;
            15'd11695: log10_cal = 16'b0000010000111011;
            15'd11696: log10_cal = 16'b0000010000111011;
            15'd11697: log10_cal = 16'b0000010000111011;
            15'd11698: log10_cal = 16'b0000010000111011;
            15'd11699: log10_cal = 16'b0000010000111011;
            15'd11700: log10_cal = 16'b0000010000111011;
            15'd11701: log10_cal = 16'b0000010000111011;
            15'd11702: log10_cal = 16'b0000010000111011;
            15'd11703: log10_cal = 16'b0000010000111011;
            15'd11704: log10_cal = 16'b0000010000111011;
            15'd11705: log10_cal = 16'b0000010000111011;
            15'd11706: log10_cal = 16'b0000010000111011;
            15'd11707: log10_cal = 16'b0000010000111011;
            15'd11708: log10_cal = 16'b0000010000111011;
            15'd11709: log10_cal = 16'b0000010000111011;
            15'd11710: log10_cal = 16'b0000010000111011;
            15'd11711: log10_cal = 16'b0000010000111011;
            15'd11712: log10_cal = 16'b0000010000111011;
            15'd11713: log10_cal = 16'b0000010000111011;
            15'd11714: log10_cal = 16'b0000010000111011;
            15'd11715: log10_cal = 16'b0000010000111011;
            15'd11716: log10_cal = 16'b0000010000111011;
            15'd11717: log10_cal = 16'b0000010000111011;
            15'd11718: log10_cal = 16'b0000010000111011;
            15'd11719: log10_cal = 16'b0000010000111011;
            15'd11720: log10_cal = 16'b0000010000111100;
            15'd11721: log10_cal = 16'b0000010000111100;
            15'd11722: log10_cal = 16'b0000010000111100;
            15'd11723: log10_cal = 16'b0000010000111100;
            15'd11724: log10_cal = 16'b0000010000111100;
            15'd11725: log10_cal = 16'b0000010000111100;
            15'd11726: log10_cal = 16'b0000010000111100;
            15'd11727: log10_cal = 16'b0000010000111100;
            15'd11728: log10_cal = 16'b0000010000111100;
            15'd11729: log10_cal = 16'b0000010000111100;
            15'd11730: log10_cal = 16'b0000010000111100;
            15'd11731: log10_cal = 16'b0000010000111100;
            15'd11732: log10_cal = 16'b0000010000111100;
            15'd11733: log10_cal = 16'b0000010000111100;
            15'd11734: log10_cal = 16'b0000010000111100;
            15'd11735: log10_cal = 16'b0000010000111100;
            15'd11736: log10_cal = 16'b0000010000111100;
            15'd11737: log10_cal = 16'b0000010000111100;
            15'd11738: log10_cal = 16'b0000010000111100;
            15'd11739: log10_cal = 16'b0000010000111100;
            15'd11740: log10_cal = 16'b0000010000111100;
            15'd11741: log10_cal = 16'b0000010000111100;
            15'd11742: log10_cal = 16'b0000010000111100;
            15'd11743: log10_cal = 16'b0000010000111100;
            15'd11744: log10_cal = 16'b0000010000111100;
            15'd11745: log10_cal = 16'b0000010000111100;
            15'd11746: log10_cal = 16'b0000010000111101;
            15'd11747: log10_cal = 16'b0000010000111101;
            15'd11748: log10_cal = 16'b0000010000111101;
            15'd11749: log10_cal = 16'b0000010000111101;
            15'd11750: log10_cal = 16'b0000010000111101;
            15'd11751: log10_cal = 16'b0000010000111101;
            15'd11752: log10_cal = 16'b0000010000111101;
            15'd11753: log10_cal = 16'b0000010000111101;
            15'd11754: log10_cal = 16'b0000010000111101;
            15'd11755: log10_cal = 16'b0000010000111101;
            15'd11756: log10_cal = 16'b0000010000111101;
            15'd11757: log10_cal = 16'b0000010000111101;
            15'd11758: log10_cal = 16'b0000010000111101;
            15'd11759: log10_cal = 16'b0000010000111101;
            15'd11760: log10_cal = 16'b0000010000111101;
            15'd11761: log10_cal = 16'b0000010000111101;
            15'd11762: log10_cal = 16'b0000010000111101;
            15'd11763: log10_cal = 16'b0000010000111101;
            15'd11764: log10_cal = 16'b0000010000111101;
            15'd11765: log10_cal = 16'b0000010000111101;
            15'd11766: log10_cal = 16'b0000010000111101;
            15'd11767: log10_cal = 16'b0000010000111101;
            15'd11768: log10_cal = 16'b0000010000111101;
            15'd11769: log10_cal = 16'b0000010000111101;
            15'd11770: log10_cal = 16'b0000010000111101;
            15'd11771: log10_cal = 16'b0000010000111101;
            15'd11772: log10_cal = 16'b0000010000111110;
            15'd11773: log10_cal = 16'b0000010000111110;
            15'd11774: log10_cal = 16'b0000010000111110;
            15'd11775: log10_cal = 16'b0000010000111110;
            15'd11776: log10_cal = 16'b0000010000111110;
            15'd11777: log10_cal = 16'b0000010000111110;
            15'd11778: log10_cal = 16'b0000010000111110;
            15'd11779: log10_cal = 16'b0000010000111110;
            15'd11780: log10_cal = 16'b0000010000111110;
            15'd11781: log10_cal = 16'b0000010000111110;
            15'd11782: log10_cal = 16'b0000010000111110;
            15'd11783: log10_cal = 16'b0000010000111110;
            15'd11784: log10_cal = 16'b0000010000111110;
            15'd11785: log10_cal = 16'b0000010000111110;
            15'd11786: log10_cal = 16'b0000010000111110;
            15'd11787: log10_cal = 16'b0000010000111110;
            15'd11788: log10_cal = 16'b0000010000111110;
            15'd11789: log10_cal = 16'b0000010000111110;
            15'd11790: log10_cal = 16'b0000010000111110;
            15'd11791: log10_cal = 16'b0000010000111110;
            15'd11792: log10_cal = 16'b0000010000111110;
            15'd11793: log10_cal = 16'b0000010000111110;
            15'd11794: log10_cal = 16'b0000010000111110;
            15'd11795: log10_cal = 16'b0000010000111110;
            15'd11796: log10_cal = 16'b0000010000111110;
            15'd11797: log10_cal = 16'b0000010000111110;
            15'd11798: log10_cal = 16'b0000010000111110;
            15'd11799: log10_cal = 16'b0000010000111111;
            15'd11800: log10_cal = 16'b0000010000111111;
            15'd11801: log10_cal = 16'b0000010000111111;
            15'd11802: log10_cal = 16'b0000010000111111;
            15'd11803: log10_cal = 16'b0000010000111111;
            15'd11804: log10_cal = 16'b0000010000111111;
            15'd11805: log10_cal = 16'b0000010000111111;
            15'd11806: log10_cal = 16'b0000010000111111;
            15'd11807: log10_cal = 16'b0000010000111111;
            15'd11808: log10_cal = 16'b0000010000111111;
            15'd11809: log10_cal = 16'b0000010000111111;
            15'd11810: log10_cal = 16'b0000010000111111;
            15'd11811: log10_cal = 16'b0000010000111111;
            15'd11812: log10_cal = 16'b0000010000111111;
            15'd11813: log10_cal = 16'b0000010000111111;
            15'd11814: log10_cal = 16'b0000010000111111;
            15'd11815: log10_cal = 16'b0000010000111111;
            15'd11816: log10_cal = 16'b0000010000111111;
            15'd11817: log10_cal = 16'b0000010000111111;
            15'd11818: log10_cal = 16'b0000010000111111;
            15'd11819: log10_cal = 16'b0000010000111111;
            15'd11820: log10_cal = 16'b0000010000111111;
            15'd11821: log10_cal = 16'b0000010000111111;
            15'd11822: log10_cal = 16'b0000010000111111;
            15'd11823: log10_cal = 16'b0000010000111111;
            15'd11824: log10_cal = 16'b0000010000111111;
            15'd11825: log10_cal = 16'b0000010001000000;
            15'd11826: log10_cal = 16'b0000010001000000;
            15'd11827: log10_cal = 16'b0000010001000000;
            15'd11828: log10_cal = 16'b0000010001000000;
            15'd11829: log10_cal = 16'b0000010001000000;
            15'd11830: log10_cal = 16'b0000010001000000;
            15'd11831: log10_cal = 16'b0000010001000000;
            15'd11832: log10_cal = 16'b0000010001000000;
            15'd11833: log10_cal = 16'b0000010001000000;
            15'd11834: log10_cal = 16'b0000010001000000;
            15'd11835: log10_cal = 16'b0000010001000000;
            15'd11836: log10_cal = 16'b0000010001000000;
            15'd11837: log10_cal = 16'b0000010001000000;
            15'd11838: log10_cal = 16'b0000010001000000;
            15'd11839: log10_cal = 16'b0000010001000000;
            15'd11840: log10_cal = 16'b0000010001000000;
            15'd11841: log10_cal = 16'b0000010001000000;
            15'd11842: log10_cal = 16'b0000010001000000;
            15'd11843: log10_cal = 16'b0000010001000000;
            15'd11844: log10_cal = 16'b0000010001000000;
            15'd11845: log10_cal = 16'b0000010001000000;
            15'd11846: log10_cal = 16'b0000010001000000;
            15'd11847: log10_cal = 16'b0000010001000000;
            15'd11848: log10_cal = 16'b0000010001000000;
            15'd11849: log10_cal = 16'b0000010001000000;
            15'd11850: log10_cal = 16'b0000010001000000;
            15'd11851: log10_cal = 16'b0000010001000000;
            15'd11852: log10_cal = 16'b0000010001000001;
            15'd11853: log10_cal = 16'b0000010001000001;
            15'd11854: log10_cal = 16'b0000010001000001;
            15'd11855: log10_cal = 16'b0000010001000001;
            15'd11856: log10_cal = 16'b0000010001000001;
            15'd11857: log10_cal = 16'b0000010001000001;
            15'd11858: log10_cal = 16'b0000010001000001;
            15'd11859: log10_cal = 16'b0000010001000001;
            15'd11860: log10_cal = 16'b0000010001000001;
            15'd11861: log10_cal = 16'b0000010001000001;
            15'd11862: log10_cal = 16'b0000010001000001;
            15'd11863: log10_cal = 16'b0000010001000001;
            15'd11864: log10_cal = 16'b0000010001000001;
            15'd11865: log10_cal = 16'b0000010001000001;
            15'd11866: log10_cal = 16'b0000010001000001;
            15'd11867: log10_cal = 16'b0000010001000001;
            15'd11868: log10_cal = 16'b0000010001000001;
            15'd11869: log10_cal = 16'b0000010001000001;
            15'd11870: log10_cal = 16'b0000010001000001;
            15'd11871: log10_cal = 16'b0000010001000001;
            15'd11872: log10_cal = 16'b0000010001000001;
            15'd11873: log10_cal = 16'b0000010001000001;
            15'd11874: log10_cal = 16'b0000010001000001;
            15'd11875: log10_cal = 16'b0000010001000001;
            15'd11876: log10_cal = 16'b0000010001000001;
            15'd11877: log10_cal = 16'b0000010001000001;
            15'd11878: log10_cal = 16'b0000010001000001;
            15'd11879: log10_cal = 16'b0000010001000010;
            15'd11880: log10_cal = 16'b0000010001000010;
            15'd11881: log10_cal = 16'b0000010001000010;
            15'd11882: log10_cal = 16'b0000010001000010;
            15'd11883: log10_cal = 16'b0000010001000010;
            15'd11884: log10_cal = 16'b0000010001000010;
            15'd11885: log10_cal = 16'b0000010001000010;
            15'd11886: log10_cal = 16'b0000010001000010;
            15'd11887: log10_cal = 16'b0000010001000010;
            15'd11888: log10_cal = 16'b0000010001000010;
            15'd11889: log10_cal = 16'b0000010001000010;
            15'd11890: log10_cal = 16'b0000010001000010;
            15'd11891: log10_cal = 16'b0000010001000010;
            15'd11892: log10_cal = 16'b0000010001000010;
            15'd11893: log10_cal = 16'b0000010001000010;
            15'd11894: log10_cal = 16'b0000010001000010;
            15'd11895: log10_cal = 16'b0000010001000010;
            15'd11896: log10_cal = 16'b0000010001000010;
            15'd11897: log10_cal = 16'b0000010001000010;
            15'd11898: log10_cal = 16'b0000010001000010;
            15'd11899: log10_cal = 16'b0000010001000010;
            15'd11900: log10_cal = 16'b0000010001000010;
            15'd11901: log10_cal = 16'b0000010001000010;
            15'd11902: log10_cal = 16'b0000010001000010;
            15'd11903: log10_cal = 16'b0000010001000010;
            15'd11904: log10_cal = 16'b0000010001000010;
            15'd11905: log10_cal = 16'b0000010001000010;
            15'd11906: log10_cal = 16'b0000010001000011;
            15'd11907: log10_cal = 16'b0000010001000011;
            15'd11908: log10_cal = 16'b0000010001000011;
            15'd11909: log10_cal = 16'b0000010001000011;
            15'd11910: log10_cal = 16'b0000010001000011;
            15'd11911: log10_cal = 16'b0000010001000011;
            15'd11912: log10_cal = 16'b0000010001000011;
            15'd11913: log10_cal = 16'b0000010001000011;
            15'd11914: log10_cal = 16'b0000010001000011;
            15'd11915: log10_cal = 16'b0000010001000011;
            15'd11916: log10_cal = 16'b0000010001000011;
            15'd11917: log10_cal = 16'b0000010001000011;
            15'd11918: log10_cal = 16'b0000010001000011;
            15'd11919: log10_cal = 16'b0000010001000011;
            15'd11920: log10_cal = 16'b0000010001000011;
            15'd11921: log10_cal = 16'b0000010001000011;
            15'd11922: log10_cal = 16'b0000010001000011;
            15'd11923: log10_cal = 16'b0000010001000011;
            15'd11924: log10_cal = 16'b0000010001000011;
            15'd11925: log10_cal = 16'b0000010001000011;
            15'd11926: log10_cal = 16'b0000010001000011;
            15'd11927: log10_cal = 16'b0000010001000011;
            15'd11928: log10_cal = 16'b0000010001000011;
            15'd11929: log10_cal = 16'b0000010001000011;
            15'd11930: log10_cal = 16'b0000010001000011;
            15'd11931: log10_cal = 16'b0000010001000011;
            15'd11932: log10_cal = 16'b0000010001000100;
            15'd11933: log10_cal = 16'b0000010001000100;
            15'd11934: log10_cal = 16'b0000010001000100;
            15'd11935: log10_cal = 16'b0000010001000100;
            15'd11936: log10_cal = 16'b0000010001000100;
            15'd11937: log10_cal = 16'b0000010001000100;
            15'd11938: log10_cal = 16'b0000010001000100;
            15'd11939: log10_cal = 16'b0000010001000100;
            15'd11940: log10_cal = 16'b0000010001000100;
            15'd11941: log10_cal = 16'b0000010001000100;
            15'd11942: log10_cal = 16'b0000010001000100;
            15'd11943: log10_cal = 16'b0000010001000100;
            15'd11944: log10_cal = 16'b0000010001000100;
            15'd11945: log10_cal = 16'b0000010001000100;
            15'd11946: log10_cal = 16'b0000010001000100;
            15'd11947: log10_cal = 16'b0000010001000100;
            15'd11948: log10_cal = 16'b0000010001000100;
            15'd11949: log10_cal = 16'b0000010001000100;
            15'd11950: log10_cal = 16'b0000010001000100;
            15'd11951: log10_cal = 16'b0000010001000100;
            15'd11952: log10_cal = 16'b0000010001000100;
            15'd11953: log10_cal = 16'b0000010001000100;
            15'd11954: log10_cal = 16'b0000010001000100;
            15'd11955: log10_cal = 16'b0000010001000100;
            15'd11956: log10_cal = 16'b0000010001000100;
            15'd11957: log10_cal = 16'b0000010001000100;
            15'd11958: log10_cal = 16'b0000010001000100;
            15'd11959: log10_cal = 16'b0000010001000101;
            15'd11960: log10_cal = 16'b0000010001000101;
            15'd11961: log10_cal = 16'b0000010001000101;
            15'd11962: log10_cal = 16'b0000010001000101;
            15'd11963: log10_cal = 16'b0000010001000101;
            15'd11964: log10_cal = 16'b0000010001000101;
            15'd11965: log10_cal = 16'b0000010001000101;
            15'd11966: log10_cal = 16'b0000010001000101;
            15'd11967: log10_cal = 16'b0000010001000101;
            15'd11968: log10_cal = 16'b0000010001000101;
            15'd11969: log10_cal = 16'b0000010001000101;
            15'd11970: log10_cal = 16'b0000010001000101;
            15'd11971: log10_cal = 16'b0000010001000101;
            15'd11972: log10_cal = 16'b0000010001000101;
            15'd11973: log10_cal = 16'b0000010001000101;
            15'd11974: log10_cal = 16'b0000010001000101;
            15'd11975: log10_cal = 16'b0000010001000101;
            15'd11976: log10_cal = 16'b0000010001000101;
            15'd11977: log10_cal = 16'b0000010001000101;
            15'd11978: log10_cal = 16'b0000010001000101;
            15'd11979: log10_cal = 16'b0000010001000101;
            15'd11980: log10_cal = 16'b0000010001000101;
            15'd11981: log10_cal = 16'b0000010001000101;
            15'd11982: log10_cal = 16'b0000010001000101;
            15'd11983: log10_cal = 16'b0000010001000101;
            15'd11984: log10_cal = 16'b0000010001000101;
            15'd11985: log10_cal = 16'b0000010001000101;
            15'd11986: log10_cal = 16'b0000010001000110;
            15'd11987: log10_cal = 16'b0000010001000110;
            15'd11988: log10_cal = 16'b0000010001000110;
            15'd11989: log10_cal = 16'b0000010001000110;
            15'd11990: log10_cal = 16'b0000010001000110;
            15'd11991: log10_cal = 16'b0000010001000110;
            15'd11992: log10_cal = 16'b0000010001000110;
            15'd11993: log10_cal = 16'b0000010001000110;
            15'd11994: log10_cal = 16'b0000010001000110;
            15'd11995: log10_cal = 16'b0000010001000110;
            15'd11996: log10_cal = 16'b0000010001000110;
            15'd11997: log10_cal = 16'b0000010001000110;
            15'd11998: log10_cal = 16'b0000010001000110;
            15'd11999: log10_cal = 16'b0000010001000110;
            15'd12000: log10_cal = 16'b0000010001000110;
            15'd12001: log10_cal = 16'b0000010001000110;
            15'd12002: log10_cal = 16'b0000010001000110;
            15'd12003: log10_cal = 16'b0000010001000110;
            15'd12004: log10_cal = 16'b0000010001000110;
            15'd12005: log10_cal = 16'b0000010001000110;
            15'd12006: log10_cal = 16'b0000010001000110;
            15'd12007: log10_cal = 16'b0000010001000110;
            15'd12008: log10_cal = 16'b0000010001000110;
            15'd12009: log10_cal = 16'b0000010001000110;
            15'd12010: log10_cal = 16'b0000010001000110;
            15'd12011: log10_cal = 16'b0000010001000110;
            15'd12012: log10_cal = 16'b0000010001000110;
            15'd12013: log10_cal = 16'b0000010001000111;
            15'd12014: log10_cal = 16'b0000010001000111;
            15'd12015: log10_cal = 16'b0000010001000111;
            15'd12016: log10_cal = 16'b0000010001000111;
            15'd12017: log10_cal = 16'b0000010001000111;
            15'd12018: log10_cal = 16'b0000010001000111;
            15'd12019: log10_cal = 16'b0000010001000111;
            15'd12020: log10_cal = 16'b0000010001000111;
            15'd12021: log10_cal = 16'b0000010001000111;
            15'd12022: log10_cal = 16'b0000010001000111;
            15'd12023: log10_cal = 16'b0000010001000111;
            15'd12024: log10_cal = 16'b0000010001000111;
            15'd12025: log10_cal = 16'b0000010001000111;
            15'd12026: log10_cal = 16'b0000010001000111;
            15'd12027: log10_cal = 16'b0000010001000111;
            15'd12028: log10_cal = 16'b0000010001000111;
            15'd12029: log10_cal = 16'b0000010001000111;
            15'd12030: log10_cal = 16'b0000010001000111;
            15'd12031: log10_cal = 16'b0000010001000111;
            15'd12032: log10_cal = 16'b0000010001000111;
            15'd12033: log10_cal = 16'b0000010001000111;
            15'd12034: log10_cal = 16'b0000010001000111;
            15'd12035: log10_cal = 16'b0000010001000111;
            15'd12036: log10_cal = 16'b0000010001000111;
            15'd12037: log10_cal = 16'b0000010001000111;
            15'd12038: log10_cal = 16'b0000010001000111;
            15'd12039: log10_cal = 16'b0000010001000111;
            15'd12040: log10_cal = 16'b0000010001001000;
            15'd12041: log10_cal = 16'b0000010001001000;
            15'd12042: log10_cal = 16'b0000010001001000;
            15'd12043: log10_cal = 16'b0000010001001000;
            15'd12044: log10_cal = 16'b0000010001001000;
            15'd12045: log10_cal = 16'b0000010001001000;
            15'd12046: log10_cal = 16'b0000010001001000;
            15'd12047: log10_cal = 16'b0000010001001000;
            15'd12048: log10_cal = 16'b0000010001001000;
            15'd12049: log10_cal = 16'b0000010001001000;
            15'd12050: log10_cal = 16'b0000010001001000;
            15'd12051: log10_cal = 16'b0000010001001000;
            15'd12052: log10_cal = 16'b0000010001001000;
            15'd12053: log10_cal = 16'b0000010001001000;
            15'd12054: log10_cal = 16'b0000010001001000;
            15'd12055: log10_cal = 16'b0000010001001000;
            15'd12056: log10_cal = 16'b0000010001001000;
            15'd12057: log10_cal = 16'b0000010001001000;
            15'd12058: log10_cal = 16'b0000010001001000;
            15'd12059: log10_cal = 16'b0000010001001000;
            15'd12060: log10_cal = 16'b0000010001001000;
            15'd12061: log10_cal = 16'b0000010001001000;
            15'd12062: log10_cal = 16'b0000010001001000;
            15'd12063: log10_cal = 16'b0000010001001000;
            15'd12064: log10_cal = 16'b0000010001001000;
            15'd12065: log10_cal = 16'b0000010001001000;
            15'd12066: log10_cal = 16'b0000010001001000;
            15'd12067: log10_cal = 16'b0000010001001001;
            15'd12068: log10_cal = 16'b0000010001001001;
            15'd12069: log10_cal = 16'b0000010001001001;
            15'd12070: log10_cal = 16'b0000010001001001;
            15'd12071: log10_cal = 16'b0000010001001001;
            15'd12072: log10_cal = 16'b0000010001001001;
            15'd12073: log10_cal = 16'b0000010001001001;
            15'd12074: log10_cal = 16'b0000010001001001;
            15'd12075: log10_cal = 16'b0000010001001001;
            15'd12076: log10_cal = 16'b0000010001001001;
            15'd12077: log10_cal = 16'b0000010001001001;
            15'd12078: log10_cal = 16'b0000010001001001;
            15'd12079: log10_cal = 16'b0000010001001001;
            15'd12080: log10_cal = 16'b0000010001001001;
            15'd12081: log10_cal = 16'b0000010001001001;
            15'd12082: log10_cal = 16'b0000010001001001;
            15'd12083: log10_cal = 16'b0000010001001001;
            15'd12084: log10_cal = 16'b0000010001001001;
            15'd12085: log10_cal = 16'b0000010001001001;
            15'd12086: log10_cal = 16'b0000010001001001;
            15'd12087: log10_cal = 16'b0000010001001001;
            15'd12088: log10_cal = 16'b0000010001001001;
            15'd12089: log10_cal = 16'b0000010001001001;
            15'd12090: log10_cal = 16'b0000010001001001;
            15'd12091: log10_cal = 16'b0000010001001001;
            15'd12092: log10_cal = 16'b0000010001001001;
            15'd12093: log10_cal = 16'b0000010001001001;
            15'd12094: log10_cal = 16'b0000010001001010;
            15'd12095: log10_cal = 16'b0000010001001010;
            15'd12096: log10_cal = 16'b0000010001001010;
            15'd12097: log10_cal = 16'b0000010001001010;
            15'd12098: log10_cal = 16'b0000010001001010;
            15'd12099: log10_cal = 16'b0000010001001010;
            15'd12100: log10_cal = 16'b0000010001001010;
            15'd12101: log10_cal = 16'b0000010001001010;
            15'd12102: log10_cal = 16'b0000010001001010;
            15'd12103: log10_cal = 16'b0000010001001010;
            15'd12104: log10_cal = 16'b0000010001001010;
            15'd12105: log10_cal = 16'b0000010001001010;
            15'd12106: log10_cal = 16'b0000010001001010;
            15'd12107: log10_cal = 16'b0000010001001010;
            15'd12108: log10_cal = 16'b0000010001001010;
            15'd12109: log10_cal = 16'b0000010001001010;
            15'd12110: log10_cal = 16'b0000010001001010;
            15'd12111: log10_cal = 16'b0000010001001010;
            15'd12112: log10_cal = 16'b0000010001001010;
            15'd12113: log10_cal = 16'b0000010001001010;
            15'd12114: log10_cal = 16'b0000010001001010;
            15'd12115: log10_cal = 16'b0000010001001010;
            15'd12116: log10_cal = 16'b0000010001001010;
            15'd12117: log10_cal = 16'b0000010001001010;
            15'd12118: log10_cal = 16'b0000010001001010;
            15'd12119: log10_cal = 16'b0000010001001010;
            15'd12120: log10_cal = 16'b0000010001001010;
            15'd12121: log10_cal = 16'b0000010001001010;
            15'd12122: log10_cal = 16'b0000010001001011;
            15'd12123: log10_cal = 16'b0000010001001011;
            15'd12124: log10_cal = 16'b0000010001001011;
            15'd12125: log10_cal = 16'b0000010001001011;
            15'd12126: log10_cal = 16'b0000010001001011;
            15'd12127: log10_cal = 16'b0000010001001011;
            15'd12128: log10_cal = 16'b0000010001001011;
            15'd12129: log10_cal = 16'b0000010001001011;
            15'd12130: log10_cal = 16'b0000010001001011;
            15'd12131: log10_cal = 16'b0000010001001011;
            15'd12132: log10_cal = 16'b0000010001001011;
            15'd12133: log10_cal = 16'b0000010001001011;
            15'd12134: log10_cal = 16'b0000010001001011;
            15'd12135: log10_cal = 16'b0000010001001011;
            15'd12136: log10_cal = 16'b0000010001001011;
            15'd12137: log10_cal = 16'b0000010001001011;
            15'd12138: log10_cal = 16'b0000010001001011;
            15'd12139: log10_cal = 16'b0000010001001011;
            15'd12140: log10_cal = 16'b0000010001001011;
            15'd12141: log10_cal = 16'b0000010001001011;
            15'd12142: log10_cal = 16'b0000010001001011;
            15'd12143: log10_cal = 16'b0000010001001011;
            15'd12144: log10_cal = 16'b0000010001001011;
            15'd12145: log10_cal = 16'b0000010001001011;
            15'd12146: log10_cal = 16'b0000010001001011;
            15'd12147: log10_cal = 16'b0000010001001011;
            15'd12148: log10_cal = 16'b0000010001001011;
            15'd12149: log10_cal = 16'b0000010001001100;
            15'd12150: log10_cal = 16'b0000010001001100;
            15'd12151: log10_cal = 16'b0000010001001100;
            15'd12152: log10_cal = 16'b0000010001001100;
            15'd12153: log10_cal = 16'b0000010001001100;
            15'd12154: log10_cal = 16'b0000010001001100;
            15'd12155: log10_cal = 16'b0000010001001100;
            15'd12156: log10_cal = 16'b0000010001001100;
            15'd12157: log10_cal = 16'b0000010001001100;
            15'd12158: log10_cal = 16'b0000010001001100;
            15'd12159: log10_cal = 16'b0000010001001100;
            15'd12160: log10_cal = 16'b0000010001001100;
            15'd12161: log10_cal = 16'b0000010001001100;
            15'd12162: log10_cal = 16'b0000010001001100;
            15'd12163: log10_cal = 16'b0000010001001100;
            15'd12164: log10_cal = 16'b0000010001001100;
            15'd12165: log10_cal = 16'b0000010001001100;
            15'd12166: log10_cal = 16'b0000010001001100;
            15'd12167: log10_cal = 16'b0000010001001100;
            15'd12168: log10_cal = 16'b0000010001001100;
            15'd12169: log10_cal = 16'b0000010001001100;
            15'd12170: log10_cal = 16'b0000010001001100;
            15'd12171: log10_cal = 16'b0000010001001100;
            15'd12172: log10_cal = 16'b0000010001001100;
            15'd12173: log10_cal = 16'b0000010001001100;
            15'd12174: log10_cal = 16'b0000010001001100;
            15'd12175: log10_cal = 16'b0000010001001100;
            15'd12176: log10_cal = 16'b0000010001001101;
            15'd12177: log10_cal = 16'b0000010001001101;
            15'd12178: log10_cal = 16'b0000010001001101;
            15'd12179: log10_cal = 16'b0000010001001101;
            15'd12180: log10_cal = 16'b0000010001001101;
            15'd12181: log10_cal = 16'b0000010001001101;
            15'd12182: log10_cal = 16'b0000010001001101;
            15'd12183: log10_cal = 16'b0000010001001101;
            15'd12184: log10_cal = 16'b0000010001001101;
            15'd12185: log10_cal = 16'b0000010001001101;
            15'd12186: log10_cal = 16'b0000010001001101;
            15'd12187: log10_cal = 16'b0000010001001101;
            15'd12188: log10_cal = 16'b0000010001001101;
            15'd12189: log10_cal = 16'b0000010001001101;
            15'd12190: log10_cal = 16'b0000010001001101;
            15'd12191: log10_cal = 16'b0000010001001101;
            15'd12192: log10_cal = 16'b0000010001001101;
            15'd12193: log10_cal = 16'b0000010001001101;
            15'd12194: log10_cal = 16'b0000010001001101;
            15'd12195: log10_cal = 16'b0000010001001101;
            15'd12196: log10_cal = 16'b0000010001001101;
            15'd12197: log10_cal = 16'b0000010001001101;
            15'd12198: log10_cal = 16'b0000010001001101;
            15'd12199: log10_cal = 16'b0000010001001101;
            15'd12200: log10_cal = 16'b0000010001001101;
            15'd12201: log10_cal = 16'b0000010001001101;
            15'd12202: log10_cal = 16'b0000010001001101;
            15'd12203: log10_cal = 16'b0000010001001101;
            15'd12204: log10_cal = 16'b0000010001001110;
            15'd12205: log10_cal = 16'b0000010001001110;
            15'd12206: log10_cal = 16'b0000010001001110;
            15'd12207: log10_cal = 16'b0000010001001110;
            15'd12208: log10_cal = 16'b0000010001001110;
            15'd12209: log10_cal = 16'b0000010001001110;
            15'd12210: log10_cal = 16'b0000010001001110;
            15'd12211: log10_cal = 16'b0000010001001110;
            15'd12212: log10_cal = 16'b0000010001001110;
            15'd12213: log10_cal = 16'b0000010001001110;
            15'd12214: log10_cal = 16'b0000010001001110;
            15'd12215: log10_cal = 16'b0000010001001110;
            15'd12216: log10_cal = 16'b0000010001001110;
            15'd12217: log10_cal = 16'b0000010001001110;
            15'd12218: log10_cal = 16'b0000010001001110;
            15'd12219: log10_cal = 16'b0000010001001110;
            15'd12220: log10_cal = 16'b0000010001001110;
            15'd12221: log10_cal = 16'b0000010001001110;
            15'd12222: log10_cal = 16'b0000010001001110;
            15'd12223: log10_cal = 16'b0000010001001110;
            15'd12224: log10_cal = 16'b0000010001001110;
            15'd12225: log10_cal = 16'b0000010001001110;
            15'd12226: log10_cal = 16'b0000010001001110;
            15'd12227: log10_cal = 16'b0000010001001110;
            15'd12228: log10_cal = 16'b0000010001001110;
            15'd12229: log10_cal = 16'b0000010001001110;
            15'd12230: log10_cal = 16'b0000010001001110;
            15'd12231: log10_cal = 16'b0000010001001111;
            15'd12232: log10_cal = 16'b0000010001001111;
            15'd12233: log10_cal = 16'b0000010001001111;
            15'd12234: log10_cal = 16'b0000010001001111;
            15'd12235: log10_cal = 16'b0000010001001111;
            15'd12236: log10_cal = 16'b0000010001001111;
            15'd12237: log10_cal = 16'b0000010001001111;
            15'd12238: log10_cal = 16'b0000010001001111;
            15'd12239: log10_cal = 16'b0000010001001111;
            15'd12240: log10_cal = 16'b0000010001001111;
            15'd12241: log10_cal = 16'b0000010001001111;
            15'd12242: log10_cal = 16'b0000010001001111;
            15'd12243: log10_cal = 16'b0000010001001111;
            15'd12244: log10_cal = 16'b0000010001001111;
            15'd12245: log10_cal = 16'b0000010001001111;
            15'd12246: log10_cal = 16'b0000010001001111;
            15'd12247: log10_cal = 16'b0000010001001111;
            15'd12248: log10_cal = 16'b0000010001001111;
            15'd12249: log10_cal = 16'b0000010001001111;
            15'd12250: log10_cal = 16'b0000010001001111;
            15'd12251: log10_cal = 16'b0000010001001111;
            15'd12252: log10_cal = 16'b0000010001001111;
            15'd12253: log10_cal = 16'b0000010001001111;
            15'd12254: log10_cal = 16'b0000010001001111;
            15'd12255: log10_cal = 16'b0000010001001111;
            15'd12256: log10_cal = 16'b0000010001001111;
            15'd12257: log10_cal = 16'b0000010001001111;
            15'd12258: log10_cal = 16'b0000010001001111;
            15'd12259: log10_cal = 16'b0000010001010000;
            15'd12260: log10_cal = 16'b0000010001010000;
            15'd12261: log10_cal = 16'b0000010001010000;
            15'd12262: log10_cal = 16'b0000010001010000;
            15'd12263: log10_cal = 16'b0000010001010000;
            15'd12264: log10_cal = 16'b0000010001010000;
            15'd12265: log10_cal = 16'b0000010001010000;
            15'd12266: log10_cal = 16'b0000010001010000;
            15'd12267: log10_cal = 16'b0000010001010000;
            15'd12268: log10_cal = 16'b0000010001010000;
            15'd12269: log10_cal = 16'b0000010001010000;
            15'd12270: log10_cal = 16'b0000010001010000;
            15'd12271: log10_cal = 16'b0000010001010000;
            15'd12272: log10_cal = 16'b0000010001010000;
            15'd12273: log10_cal = 16'b0000010001010000;
            15'd12274: log10_cal = 16'b0000010001010000;
            15'd12275: log10_cal = 16'b0000010001010000;
            15'd12276: log10_cal = 16'b0000010001010000;
            15'd12277: log10_cal = 16'b0000010001010000;
            15'd12278: log10_cal = 16'b0000010001010000;
            15'd12279: log10_cal = 16'b0000010001010000;
            15'd12280: log10_cal = 16'b0000010001010000;
            15'd12281: log10_cal = 16'b0000010001010000;
            15'd12282: log10_cal = 16'b0000010001010000;
            15'd12283: log10_cal = 16'b0000010001010000;
            15'd12284: log10_cal = 16'b0000010001010000;
            15'd12285: log10_cal = 16'b0000010001010000;
            15'd12286: log10_cal = 16'b0000010001010001;
            15'd12287: log10_cal = 16'b0000010001010001;
            15'd12288: log10_cal = 16'b0000010001010001;
            15'd12289: log10_cal = 16'b0000010001010001;
            15'd12290: log10_cal = 16'b0000010001010001;
            15'd12291: log10_cal = 16'b0000010001010001;
            15'd12292: log10_cal = 16'b0000010001010001;
            15'd12293: log10_cal = 16'b0000010001010001;
            15'd12294: log10_cal = 16'b0000010001010001;
            15'd12295: log10_cal = 16'b0000010001010001;
            15'd12296: log10_cal = 16'b0000010001010001;
            15'd12297: log10_cal = 16'b0000010001010001;
            15'd12298: log10_cal = 16'b0000010001010001;
            15'd12299: log10_cal = 16'b0000010001010001;
            15'd12300: log10_cal = 16'b0000010001010001;
            15'd12301: log10_cal = 16'b0000010001010001;
            15'd12302: log10_cal = 16'b0000010001010001;
            15'd12303: log10_cal = 16'b0000010001010001;
            15'd12304: log10_cal = 16'b0000010001010001;
            15'd12305: log10_cal = 16'b0000010001010001;
            15'd12306: log10_cal = 16'b0000010001010001;
            15'd12307: log10_cal = 16'b0000010001010001;
            15'd12308: log10_cal = 16'b0000010001010001;
            15'd12309: log10_cal = 16'b0000010001010001;
            15'd12310: log10_cal = 16'b0000010001010001;
            15'd12311: log10_cal = 16'b0000010001010001;
            15'd12312: log10_cal = 16'b0000010001010001;
            15'd12313: log10_cal = 16'b0000010001010001;
            15'd12314: log10_cal = 16'b0000010001010010;
            15'd12315: log10_cal = 16'b0000010001010010;
            15'd12316: log10_cal = 16'b0000010001010010;
            15'd12317: log10_cal = 16'b0000010001010010;
            15'd12318: log10_cal = 16'b0000010001010010;
            15'd12319: log10_cal = 16'b0000010001010010;
            15'd12320: log10_cal = 16'b0000010001010010;
            15'd12321: log10_cal = 16'b0000010001010010;
            15'd12322: log10_cal = 16'b0000010001010010;
            15'd12323: log10_cal = 16'b0000010001010010;
            15'd12324: log10_cal = 16'b0000010001010010;
            15'd12325: log10_cal = 16'b0000010001010010;
            15'd12326: log10_cal = 16'b0000010001010010;
            15'd12327: log10_cal = 16'b0000010001010010;
            15'd12328: log10_cal = 16'b0000010001010010;
            15'd12329: log10_cal = 16'b0000010001010010;
            15'd12330: log10_cal = 16'b0000010001010010;
            15'd12331: log10_cal = 16'b0000010001010010;
            15'd12332: log10_cal = 16'b0000010001010010;
            15'd12333: log10_cal = 16'b0000010001010010;
            15'd12334: log10_cal = 16'b0000010001010010;
            15'd12335: log10_cal = 16'b0000010001010010;
            15'd12336: log10_cal = 16'b0000010001010010;
            15'd12337: log10_cal = 16'b0000010001010010;
            15'd12338: log10_cal = 16'b0000010001010010;
            15'd12339: log10_cal = 16'b0000010001010010;
            15'd12340: log10_cal = 16'b0000010001010010;
            15'd12341: log10_cal = 16'b0000010001010010;
            15'd12342: log10_cal = 16'b0000010001010011;
            15'd12343: log10_cal = 16'b0000010001010011;
            15'd12344: log10_cal = 16'b0000010001010011;
            15'd12345: log10_cal = 16'b0000010001010011;
            15'd12346: log10_cal = 16'b0000010001010011;
            15'd12347: log10_cal = 16'b0000010001010011;
            15'd12348: log10_cal = 16'b0000010001010011;
            15'd12349: log10_cal = 16'b0000010001010011;
            15'd12350: log10_cal = 16'b0000010001010011;
            15'd12351: log10_cal = 16'b0000010001010011;
            15'd12352: log10_cal = 16'b0000010001010011;
            15'd12353: log10_cal = 16'b0000010001010011;
            15'd12354: log10_cal = 16'b0000010001010011;
            15'd12355: log10_cal = 16'b0000010001010011;
            15'd12356: log10_cal = 16'b0000010001010011;
            15'd12357: log10_cal = 16'b0000010001010011;
            15'd12358: log10_cal = 16'b0000010001010011;
            15'd12359: log10_cal = 16'b0000010001010011;
            15'd12360: log10_cal = 16'b0000010001010011;
            15'd12361: log10_cal = 16'b0000010001010011;
            15'd12362: log10_cal = 16'b0000010001010011;
            15'd12363: log10_cal = 16'b0000010001010011;
            15'd12364: log10_cal = 16'b0000010001010011;
            15'd12365: log10_cal = 16'b0000010001010011;
            15'd12366: log10_cal = 16'b0000010001010011;
            15'd12367: log10_cal = 16'b0000010001010011;
            15'd12368: log10_cal = 16'b0000010001010011;
            15'd12369: log10_cal = 16'b0000010001010100;
            15'd12370: log10_cal = 16'b0000010001010100;
            15'd12371: log10_cal = 16'b0000010001010100;
            15'd12372: log10_cal = 16'b0000010001010100;
            15'd12373: log10_cal = 16'b0000010001010100;
            15'd12374: log10_cal = 16'b0000010001010100;
            15'd12375: log10_cal = 16'b0000010001010100;
            15'd12376: log10_cal = 16'b0000010001010100;
            15'd12377: log10_cal = 16'b0000010001010100;
            15'd12378: log10_cal = 16'b0000010001010100;
            15'd12379: log10_cal = 16'b0000010001010100;
            15'd12380: log10_cal = 16'b0000010001010100;
            15'd12381: log10_cal = 16'b0000010001010100;
            15'd12382: log10_cal = 16'b0000010001010100;
            15'd12383: log10_cal = 16'b0000010001010100;
            15'd12384: log10_cal = 16'b0000010001010100;
            15'd12385: log10_cal = 16'b0000010001010100;
            15'd12386: log10_cal = 16'b0000010001010100;
            15'd12387: log10_cal = 16'b0000010001010100;
            15'd12388: log10_cal = 16'b0000010001010100;
            15'd12389: log10_cal = 16'b0000010001010100;
            15'd12390: log10_cal = 16'b0000010001010100;
            15'd12391: log10_cal = 16'b0000010001010100;
            15'd12392: log10_cal = 16'b0000010001010100;
            15'd12393: log10_cal = 16'b0000010001010100;
            15'd12394: log10_cal = 16'b0000010001010100;
            15'd12395: log10_cal = 16'b0000010001010100;
            15'd12396: log10_cal = 16'b0000010001010100;
            15'd12397: log10_cal = 16'b0000010001010101;
            15'd12398: log10_cal = 16'b0000010001010101;
            15'd12399: log10_cal = 16'b0000010001010101;
            15'd12400: log10_cal = 16'b0000010001010101;
            15'd12401: log10_cal = 16'b0000010001010101;
            15'd12402: log10_cal = 16'b0000010001010101;
            15'd12403: log10_cal = 16'b0000010001010101;
            15'd12404: log10_cal = 16'b0000010001010101;
            15'd12405: log10_cal = 16'b0000010001010101;
            15'd12406: log10_cal = 16'b0000010001010101;
            15'd12407: log10_cal = 16'b0000010001010101;
            15'd12408: log10_cal = 16'b0000010001010101;
            15'd12409: log10_cal = 16'b0000010001010101;
            15'd12410: log10_cal = 16'b0000010001010101;
            15'd12411: log10_cal = 16'b0000010001010101;
            15'd12412: log10_cal = 16'b0000010001010101;
            15'd12413: log10_cal = 16'b0000010001010101;
            15'd12414: log10_cal = 16'b0000010001010101;
            15'd12415: log10_cal = 16'b0000010001010101;
            15'd12416: log10_cal = 16'b0000010001010101;
            15'd12417: log10_cal = 16'b0000010001010101;
            15'd12418: log10_cal = 16'b0000010001010101;
            15'd12419: log10_cal = 16'b0000010001010101;
            15'd12420: log10_cal = 16'b0000010001010101;
            15'd12421: log10_cal = 16'b0000010001010101;
            15'd12422: log10_cal = 16'b0000010001010101;
            15'd12423: log10_cal = 16'b0000010001010101;
            15'd12424: log10_cal = 16'b0000010001010101;
            15'd12425: log10_cal = 16'b0000010001010110;
            15'd12426: log10_cal = 16'b0000010001010110;
            15'd12427: log10_cal = 16'b0000010001010110;
            15'd12428: log10_cal = 16'b0000010001010110;
            15'd12429: log10_cal = 16'b0000010001010110;
            15'd12430: log10_cal = 16'b0000010001010110;
            15'd12431: log10_cal = 16'b0000010001010110;
            15'd12432: log10_cal = 16'b0000010001010110;
            15'd12433: log10_cal = 16'b0000010001010110;
            15'd12434: log10_cal = 16'b0000010001010110;
            15'd12435: log10_cal = 16'b0000010001010110;
            15'd12436: log10_cal = 16'b0000010001010110;
            15'd12437: log10_cal = 16'b0000010001010110;
            15'd12438: log10_cal = 16'b0000010001010110;
            15'd12439: log10_cal = 16'b0000010001010110;
            15'd12440: log10_cal = 16'b0000010001010110;
            15'd12441: log10_cal = 16'b0000010001010110;
            15'd12442: log10_cal = 16'b0000010001010110;
            15'd12443: log10_cal = 16'b0000010001010110;
            15'd12444: log10_cal = 16'b0000010001010110;
            15'd12445: log10_cal = 16'b0000010001010110;
            15'd12446: log10_cal = 16'b0000010001010110;
            15'd12447: log10_cal = 16'b0000010001010110;
            15'd12448: log10_cal = 16'b0000010001010110;
            15'd12449: log10_cal = 16'b0000010001010110;
            15'd12450: log10_cal = 16'b0000010001010110;
            15'd12451: log10_cal = 16'b0000010001010110;
            15'd12452: log10_cal = 16'b0000010001010110;
            15'd12453: log10_cal = 16'b0000010001010111;
            15'd12454: log10_cal = 16'b0000010001010111;
            15'd12455: log10_cal = 16'b0000010001010111;
            15'd12456: log10_cal = 16'b0000010001010111;
            15'd12457: log10_cal = 16'b0000010001010111;
            15'd12458: log10_cal = 16'b0000010001010111;
            15'd12459: log10_cal = 16'b0000010001010111;
            15'd12460: log10_cal = 16'b0000010001010111;
            15'd12461: log10_cal = 16'b0000010001010111;
            15'd12462: log10_cal = 16'b0000010001010111;
            15'd12463: log10_cal = 16'b0000010001010111;
            15'd12464: log10_cal = 16'b0000010001010111;
            15'd12465: log10_cal = 16'b0000010001010111;
            15'd12466: log10_cal = 16'b0000010001010111;
            15'd12467: log10_cal = 16'b0000010001010111;
            15'd12468: log10_cal = 16'b0000010001010111;
            15'd12469: log10_cal = 16'b0000010001010111;
            15'd12470: log10_cal = 16'b0000010001010111;
            15'd12471: log10_cal = 16'b0000010001010111;
            15'd12472: log10_cal = 16'b0000010001010111;
            15'd12473: log10_cal = 16'b0000010001010111;
            15'd12474: log10_cal = 16'b0000010001010111;
            15'd12475: log10_cal = 16'b0000010001010111;
            15'd12476: log10_cal = 16'b0000010001010111;
            15'd12477: log10_cal = 16'b0000010001010111;
            15'd12478: log10_cal = 16'b0000010001010111;
            15'd12479: log10_cal = 16'b0000010001010111;
            15'd12480: log10_cal = 16'b0000010001010111;
            15'd12481: log10_cal = 16'b0000010001011000;
            15'd12482: log10_cal = 16'b0000010001011000;
            15'd12483: log10_cal = 16'b0000010001011000;
            15'd12484: log10_cal = 16'b0000010001011000;
            15'd12485: log10_cal = 16'b0000010001011000;
            15'd12486: log10_cal = 16'b0000010001011000;
            15'd12487: log10_cal = 16'b0000010001011000;
            15'd12488: log10_cal = 16'b0000010001011000;
            15'd12489: log10_cal = 16'b0000010001011000;
            15'd12490: log10_cal = 16'b0000010001011000;
            15'd12491: log10_cal = 16'b0000010001011000;
            15'd12492: log10_cal = 16'b0000010001011000;
            15'd12493: log10_cal = 16'b0000010001011000;
            15'd12494: log10_cal = 16'b0000010001011000;
            15'd12495: log10_cal = 16'b0000010001011000;
            15'd12496: log10_cal = 16'b0000010001011000;
            15'd12497: log10_cal = 16'b0000010001011000;
            15'd12498: log10_cal = 16'b0000010001011000;
            15'd12499: log10_cal = 16'b0000010001011000;
            15'd12500: log10_cal = 16'b0000010001011000;
            15'd12501: log10_cal = 16'b0000010001011000;
            15'd12502: log10_cal = 16'b0000010001011000;
            15'd12503: log10_cal = 16'b0000010001011000;
            15'd12504: log10_cal = 16'b0000010001011000;
            15'd12505: log10_cal = 16'b0000010001011000;
            15'd12506: log10_cal = 16'b0000010001011000;
            15'd12507: log10_cal = 16'b0000010001011000;
            15'd12508: log10_cal = 16'b0000010001011000;
            15'd12509: log10_cal = 16'b0000010001011001;
            15'd12510: log10_cal = 16'b0000010001011001;
            15'd12511: log10_cal = 16'b0000010001011001;
            15'd12512: log10_cal = 16'b0000010001011001;
            15'd12513: log10_cal = 16'b0000010001011001;
            15'd12514: log10_cal = 16'b0000010001011001;
            15'd12515: log10_cal = 16'b0000010001011001;
            15'd12516: log10_cal = 16'b0000010001011001;
            15'd12517: log10_cal = 16'b0000010001011001;
            15'd12518: log10_cal = 16'b0000010001011001;
            15'd12519: log10_cal = 16'b0000010001011001;
            15'd12520: log10_cal = 16'b0000010001011001;
            15'd12521: log10_cal = 16'b0000010001011001;
            15'd12522: log10_cal = 16'b0000010001011001;
            15'd12523: log10_cal = 16'b0000010001011001;
            15'd12524: log10_cal = 16'b0000010001011001;
            15'd12525: log10_cal = 16'b0000010001011001;
            15'd12526: log10_cal = 16'b0000010001011001;
            15'd12527: log10_cal = 16'b0000010001011001;
            15'd12528: log10_cal = 16'b0000010001011001;
            15'd12529: log10_cal = 16'b0000010001011001;
            15'd12530: log10_cal = 16'b0000010001011001;
            15'd12531: log10_cal = 16'b0000010001011001;
            15'd12532: log10_cal = 16'b0000010001011001;
            15'd12533: log10_cal = 16'b0000010001011001;
            15'd12534: log10_cal = 16'b0000010001011001;
            15'd12535: log10_cal = 16'b0000010001011001;
            15'd12536: log10_cal = 16'b0000010001011001;
            15'd12537: log10_cal = 16'b0000010001011010;
            15'd12538: log10_cal = 16'b0000010001011010;
            15'd12539: log10_cal = 16'b0000010001011010;
            15'd12540: log10_cal = 16'b0000010001011010;
            15'd12541: log10_cal = 16'b0000010001011010;
            15'd12542: log10_cal = 16'b0000010001011010;
            15'd12543: log10_cal = 16'b0000010001011010;
            15'd12544: log10_cal = 16'b0000010001011010;
            15'd12545: log10_cal = 16'b0000010001011010;
            15'd12546: log10_cal = 16'b0000010001011010;
            15'd12547: log10_cal = 16'b0000010001011010;
            15'd12548: log10_cal = 16'b0000010001011010;
            15'd12549: log10_cal = 16'b0000010001011010;
            15'd12550: log10_cal = 16'b0000010001011010;
            15'd12551: log10_cal = 16'b0000010001011010;
            15'd12552: log10_cal = 16'b0000010001011010;
            15'd12553: log10_cal = 16'b0000010001011010;
            15'd12554: log10_cal = 16'b0000010001011010;
            15'd12555: log10_cal = 16'b0000010001011010;
            15'd12556: log10_cal = 16'b0000010001011010;
            15'd12557: log10_cal = 16'b0000010001011010;
            15'd12558: log10_cal = 16'b0000010001011010;
            15'd12559: log10_cal = 16'b0000010001011010;
            15'd12560: log10_cal = 16'b0000010001011010;
            15'd12561: log10_cal = 16'b0000010001011010;
            15'd12562: log10_cal = 16'b0000010001011010;
            15'd12563: log10_cal = 16'b0000010001011010;
            15'd12564: log10_cal = 16'b0000010001011010;
            15'd12565: log10_cal = 16'b0000010001011010;
            15'd12566: log10_cal = 16'b0000010001011011;
            15'd12567: log10_cal = 16'b0000010001011011;
            15'd12568: log10_cal = 16'b0000010001011011;
            15'd12569: log10_cal = 16'b0000010001011011;
            15'd12570: log10_cal = 16'b0000010001011011;
            15'd12571: log10_cal = 16'b0000010001011011;
            15'd12572: log10_cal = 16'b0000010001011011;
            15'd12573: log10_cal = 16'b0000010001011011;
            15'd12574: log10_cal = 16'b0000010001011011;
            15'd12575: log10_cal = 16'b0000010001011011;
            15'd12576: log10_cal = 16'b0000010001011011;
            15'd12577: log10_cal = 16'b0000010001011011;
            15'd12578: log10_cal = 16'b0000010001011011;
            15'd12579: log10_cal = 16'b0000010001011011;
            15'd12580: log10_cal = 16'b0000010001011011;
            15'd12581: log10_cal = 16'b0000010001011011;
            15'd12582: log10_cal = 16'b0000010001011011;
            15'd12583: log10_cal = 16'b0000010001011011;
            15'd12584: log10_cal = 16'b0000010001011011;
            15'd12585: log10_cal = 16'b0000010001011011;
            15'd12586: log10_cal = 16'b0000010001011011;
            15'd12587: log10_cal = 16'b0000010001011011;
            15'd12588: log10_cal = 16'b0000010001011011;
            15'd12589: log10_cal = 16'b0000010001011011;
            15'd12590: log10_cal = 16'b0000010001011011;
            15'd12591: log10_cal = 16'b0000010001011011;
            15'd12592: log10_cal = 16'b0000010001011011;
            15'd12593: log10_cal = 16'b0000010001011011;
            15'd12594: log10_cal = 16'b0000010001011100;
            15'd12595: log10_cal = 16'b0000010001011100;
            15'd12596: log10_cal = 16'b0000010001011100;
            15'd12597: log10_cal = 16'b0000010001011100;
            15'd12598: log10_cal = 16'b0000010001011100;
            15'd12599: log10_cal = 16'b0000010001011100;
            15'd12600: log10_cal = 16'b0000010001011100;
            15'd12601: log10_cal = 16'b0000010001011100;
            15'd12602: log10_cal = 16'b0000010001011100;
            15'd12603: log10_cal = 16'b0000010001011100;
            15'd12604: log10_cal = 16'b0000010001011100;
            15'd12605: log10_cal = 16'b0000010001011100;
            15'd12606: log10_cal = 16'b0000010001011100;
            15'd12607: log10_cal = 16'b0000010001011100;
            15'd12608: log10_cal = 16'b0000010001011100;
            15'd12609: log10_cal = 16'b0000010001011100;
            15'd12610: log10_cal = 16'b0000010001011100;
            15'd12611: log10_cal = 16'b0000010001011100;
            15'd12612: log10_cal = 16'b0000010001011100;
            15'd12613: log10_cal = 16'b0000010001011100;
            15'd12614: log10_cal = 16'b0000010001011100;
            15'd12615: log10_cal = 16'b0000010001011100;
            15'd12616: log10_cal = 16'b0000010001011100;
            15'd12617: log10_cal = 16'b0000010001011100;
            15'd12618: log10_cal = 16'b0000010001011100;
            15'd12619: log10_cal = 16'b0000010001011100;
            15'd12620: log10_cal = 16'b0000010001011100;
            15'd12621: log10_cal = 16'b0000010001011100;
            15'd12622: log10_cal = 16'b0000010001011101;
            15'd12623: log10_cal = 16'b0000010001011101;
            15'd12624: log10_cal = 16'b0000010001011101;
            15'd12625: log10_cal = 16'b0000010001011101;
            15'd12626: log10_cal = 16'b0000010001011101;
            15'd12627: log10_cal = 16'b0000010001011101;
            15'd12628: log10_cal = 16'b0000010001011101;
            15'd12629: log10_cal = 16'b0000010001011101;
            15'd12630: log10_cal = 16'b0000010001011101;
            15'd12631: log10_cal = 16'b0000010001011101;
            15'd12632: log10_cal = 16'b0000010001011101;
            15'd12633: log10_cal = 16'b0000010001011101;
            15'd12634: log10_cal = 16'b0000010001011101;
            15'd12635: log10_cal = 16'b0000010001011101;
            15'd12636: log10_cal = 16'b0000010001011101;
            15'd12637: log10_cal = 16'b0000010001011101;
            15'd12638: log10_cal = 16'b0000010001011101;
            15'd12639: log10_cal = 16'b0000010001011101;
            15'd12640: log10_cal = 16'b0000010001011101;
            15'd12641: log10_cal = 16'b0000010001011101;
            15'd12642: log10_cal = 16'b0000010001011101;
            15'd12643: log10_cal = 16'b0000010001011101;
            15'd12644: log10_cal = 16'b0000010001011101;
            15'd12645: log10_cal = 16'b0000010001011101;
            15'd12646: log10_cal = 16'b0000010001011101;
            15'd12647: log10_cal = 16'b0000010001011101;
            15'd12648: log10_cal = 16'b0000010001011101;
            15'd12649: log10_cal = 16'b0000010001011101;
            15'd12650: log10_cal = 16'b0000010001011101;
            15'd12651: log10_cal = 16'b0000010001011110;
            15'd12652: log10_cal = 16'b0000010001011110;
            15'd12653: log10_cal = 16'b0000010001011110;
            15'd12654: log10_cal = 16'b0000010001011110;
            15'd12655: log10_cal = 16'b0000010001011110;
            15'd12656: log10_cal = 16'b0000010001011110;
            15'd12657: log10_cal = 16'b0000010001011110;
            15'd12658: log10_cal = 16'b0000010001011110;
            15'd12659: log10_cal = 16'b0000010001011110;
            15'd12660: log10_cal = 16'b0000010001011110;
            15'd12661: log10_cal = 16'b0000010001011110;
            15'd12662: log10_cal = 16'b0000010001011110;
            15'd12663: log10_cal = 16'b0000010001011110;
            15'd12664: log10_cal = 16'b0000010001011110;
            15'd12665: log10_cal = 16'b0000010001011110;
            15'd12666: log10_cal = 16'b0000010001011110;
            15'd12667: log10_cal = 16'b0000010001011110;
            15'd12668: log10_cal = 16'b0000010001011110;
            15'd12669: log10_cal = 16'b0000010001011110;
            15'd12670: log10_cal = 16'b0000010001011110;
            15'd12671: log10_cal = 16'b0000010001011110;
            15'd12672: log10_cal = 16'b0000010001011110;
            15'd12673: log10_cal = 16'b0000010001011110;
            15'd12674: log10_cal = 16'b0000010001011110;
            15'd12675: log10_cal = 16'b0000010001011110;
            15'd12676: log10_cal = 16'b0000010001011110;
            15'd12677: log10_cal = 16'b0000010001011110;
            15'd12678: log10_cal = 16'b0000010001011110;
            15'd12679: log10_cal = 16'b0000010001011111;
            15'd12680: log10_cal = 16'b0000010001011111;
            15'd12681: log10_cal = 16'b0000010001011111;
            15'd12682: log10_cal = 16'b0000010001011111;
            15'd12683: log10_cal = 16'b0000010001011111;
            15'd12684: log10_cal = 16'b0000010001011111;
            15'd12685: log10_cal = 16'b0000010001011111;
            15'd12686: log10_cal = 16'b0000010001011111;
            15'd12687: log10_cal = 16'b0000010001011111;
            15'd12688: log10_cal = 16'b0000010001011111;
            15'd12689: log10_cal = 16'b0000010001011111;
            15'd12690: log10_cal = 16'b0000010001011111;
            15'd12691: log10_cal = 16'b0000010001011111;
            15'd12692: log10_cal = 16'b0000010001011111;
            15'd12693: log10_cal = 16'b0000010001011111;
            15'd12694: log10_cal = 16'b0000010001011111;
            15'd12695: log10_cal = 16'b0000010001011111;
            15'd12696: log10_cal = 16'b0000010001011111;
            15'd12697: log10_cal = 16'b0000010001011111;
            15'd12698: log10_cal = 16'b0000010001011111;
            15'd12699: log10_cal = 16'b0000010001011111;
            15'd12700: log10_cal = 16'b0000010001011111;
            15'd12701: log10_cal = 16'b0000010001011111;
            15'd12702: log10_cal = 16'b0000010001011111;
            15'd12703: log10_cal = 16'b0000010001011111;
            15'd12704: log10_cal = 16'b0000010001011111;
            15'd12705: log10_cal = 16'b0000010001011111;
            15'd12706: log10_cal = 16'b0000010001011111;
            15'd12707: log10_cal = 16'b0000010001011111;
            15'd12708: log10_cal = 16'b0000010001100000;
            15'd12709: log10_cal = 16'b0000010001100000;
            15'd12710: log10_cal = 16'b0000010001100000;
            15'd12711: log10_cal = 16'b0000010001100000;
            15'd12712: log10_cal = 16'b0000010001100000;
            15'd12713: log10_cal = 16'b0000010001100000;
            15'd12714: log10_cal = 16'b0000010001100000;
            15'd12715: log10_cal = 16'b0000010001100000;
            15'd12716: log10_cal = 16'b0000010001100000;
            15'd12717: log10_cal = 16'b0000010001100000;
            15'd12718: log10_cal = 16'b0000010001100000;
            15'd12719: log10_cal = 16'b0000010001100000;
            15'd12720: log10_cal = 16'b0000010001100000;
            15'd12721: log10_cal = 16'b0000010001100000;
            15'd12722: log10_cal = 16'b0000010001100000;
            15'd12723: log10_cal = 16'b0000010001100000;
            15'd12724: log10_cal = 16'b0000010001100000;
            15'd12725: log10_cal = 16'b0000010001100000;
            15'd12726: log10_cal = 16'b0000010001100000;
            15'd12727: log10_cal = 16'b0000010001100000;
            15'd12728: log10_cal = 16'b0000010001100000;
            15'd12729: log10_cal = 16'b0000010001100000;
            15'd12730: log10_cal = 16'b0000010001100000;
            15'd12731: log10_cal = 16'b0000010001100000;
            15'd12732: log10_cal = 16'b0000010001100000;
            15'd12733: log10_cal = 16'b0000010001100000;
            15'd12734: log10_cal = 16'b0000010001100000;
            15'd12735: log10_cal = 16'b0000010001100000;
            15'd12736: log10_cal = 16'b0000010001100001;
            15'd12737: log10_cal = 16'b0000010001100001;
            15'd12738: log10_cal = 16'b0000010001100001;
            15'd12739: log10_cal = 16'b0000010001100001;
            15'd12740: log10_cal = 16'b0000010001100001;
            15'd12741: log10_cal = 16'b0000010001100001;
            15'd12742: log10_cal = 16'b0000010001100001;
            15'd12743: log10_cal = 16'b0000010001100001;
            15'd12744: log10_cal = 16'b0000010001100001;
            15'd12745: log10_cal = 16'b0000010001100001;
            15'd12746: log10_cal = 16'b0000010001100001;
            15'd12747: log10_cal = 16'b0000010001100001;
            15'd12748: log10_cal = 16'b0000010001100001;
            15'd12749: log10_cal = 16'b0000010001100001;
            15'd12750: log10_cal = 16'b0000010001100001;
            15'd12751: log10_cal = 16'b0000010001100001;
            15'd12752: log10_cal = 16'b0000010001100001;
            15'd12753: log10_cal = 16'b0000010001100001;
            15'd12754: log10_cal = 16'b0000010001100001;
            15'd12755: log10_cal = 16'b0000010001100001;
            15'd12756: log10_cal = 16'b0000010001100001;
            15'd12757: log10_cal = 16'b0000010001100001;
            15'd12758: log10_cal = 16'b0000010001100001;
            15'd12759: log10_cal = 16'b0000010001100001;
            15'd12760: log10_cal = 16'b0000010001100001;
            15'd12761: log10_cal = 16'b0000010001100001;
            15'd12762: log10_cal = 16'b0000010001100001;
            15'd12763: log10_cal = 16'b0000010001100001;
            15'd12764: log10_cal = 16'b0000010001100001;
            15'd12765: log10_cal = 16'b0000010001100010;
            15'd12766: log10_cal = 16'b0000010001100010;
            15'd12767: log10_cal = 16'b0000010001100010;
            15'd12768: log10_cal = 16'b0000010001100010;
            15'd12769: log10_cal = 16'b0000010001100010;
            15'd12770: log10_cal = 16'b0000010001100010;
            15'd12771: log10_cal = 16'b0000010001100010;
            15'd12772: log10_cal = 16'b0000010001100010;
            15'd12773: log10_cal = 16'b0000010001100010;
            15'd12774: log10_cal = 16'b0000010001100010;
            15'd12775: log10_cal = 16'b0000010001100010;
            15'd12776: log10_cal = 16'b0000010001100010;
            15'd12777: log10_cal = 16'b0000010001100010;
            15'd12778: log10_cal = 16'b0000010001100010;
            15'd12779: log10_cal = 16'b0000010001100010;
            15'd12780: log10_cal = 16'b0000010001100010;
            15'd12781: log10_cal = 16'b0000010001100010;
            15'd12782: log10_cal = 16'b0000010001100010;
            15'd12783: log10_cal = 16'b0000010001100010;
            15'd12784: log10_cal = 16'b0000010001100010;
            15'd12785: log10_cal = 16'b0000010001100010;
            15'd12786: log10_cal = 16'b0000010001100010;
            15'd12787: log10_cal = 16'b0000010001100010;
            15'd12788: log10_cal = 16'b0000010001100010;
            15'd12789: log10_cal = 16'b0000010001100010;
            15'd12790: log10_cal = 16'b0000010001100010;
            15'd12791: log10_cal = 16'b0000010001100010;
            15'd12792: log10_cal = 16'b0000010001100010;
            15'd12793: log10_cal = 16'b0000010001100010;
            15'd12794: log10_cal = 16'b0000010001100011;
            15'd12795: log10_cal = 16'b0000010001100011;
            15'd12796: log10_cal = 16'b0000010001100011;
            15'd12797: log10_cal = 16'b0000010001100011;
            15'd12798: log10_cal = 16'b0000010001100011;
            15'd12799: log10_cal = 16'b0000010001100011;
            15'd12800: log10_cal = 16'b0000010001100011;
            15'd12801: log10_cal = 16'b0000010001100011;
            15'd12802: log10_cal = 16'b0000010001100011;
            15'd12803: log10_cal = 16'b0000010001100011;
            15'd12804: log10_cal = 16'b0000010001100011;
            15'd12805: log10_cal = 16'b0000010001100011;
            15'd12806: log10_cal = 16'b0000010001100011;
            15'd12807: log10_cal = 16'b0000010001100011;
            15'd12808: log10_cal = 16'b0000010001100011;
            15'd12809: log10_cal = 16'b0000010001100011;
            15'd12810: log10_cal = 16'b0000010001100011;
            15'd12811: log10_cal = 16'b0000010001100011;
            15'd12812: log10_cal = 16'b0000010001100011;
            15'd12813: log10_cal = 16'b0000010001100011;
            15'd12814: log10_cal = 16'b0000010001100011;
            15'd12815: log10_cal = 16'b0000010001100011;
            15'd12816: log10_cal = 16'b0000010001100011;
            15'd12817: log10_cal = 16'b0000010001100011;
            15'd12818: log10_cal = 16'b0000010001100011;
            15'd12819: log10_cal = 16'b0000010001100011;
            15'd12820: log10_cal = 16'b0000010001100011;
            15'd12821: log10_cal = 16'b0000010001100011;
            15'd12822: log10_cal = 16'b0000010001100011;
            15'd12823: log10_cal = 16'b0000010001100100;
            15'd12824: log10_cal = 16'b0000010001100100;
            15'd12825: log10_cal = 16'b0000010001100100;
            15'd12826: log10_cal = 16'b0000010001100100;
            15'd12827: log10_cal = 16'b0000010001100100;
            15'd12828: log10_cal = 16'b0000010001100100;
            15'd12829: log10_cal = 16'b0000010001100100;
            15'd12830: log10_cal = 16'b0000010001100100;
            15'd12831: log10_cal = 16'b0000010001100100;
            15'd12832: log10_cal = 16'b0000010001100100;
            15'd12833: log10_cal = 16'b0000010001100100;
            15'd12834: log10_cal = 16'b0000010001100100;
            15'd12835: log10_cal = 16'b0000010001100100;
            15'd12836: log10_cal = 16'b0000010001100100;
            15'd12837: log10_cal = 16'b0000010001100100;
            15'd12838: log10_cal = 16'b0000010001100100;
            15'd12839: log10_cal = 16'b0000010001100100;
            15'd12840: log10_cal = 16'b0000010001100100;
            15'd12841: log10_cal = 16'b0000010001100100;
            15'd12842: log10_cal = 16'b0000010001100100;
            15'd12843: log10_cal = 16'b0000010001100100;
            15'd12844: log10_cal = 16'b0000010001100100;
            15'd12845: log10_cal = 16'b0000010001100100;
            15'd12846: log10_cal = 16'b0000010001100100;
            15'd12847: log10_cal = 16'b0000010001100100;
            15'd12848: log10_cal = 16'b0000010001100100;
            15'd12849: log10_cal = 16'b0000010001100100;
            15'd12850: log10_cal = 16'b0000010001100100;
            15'd12851: log10_cal = 16'b0000010001100101;
            15'd12852: log10_cal = 16'b0000010001100101;
            15'd12853: log10_cal = 16'b0000010001100101;
            15'd12854: log10_cal = 16'b0000010001100101;
            15'd12855: log10_cal = 16'b0000010001100101;
            15'd12856: log10_cal = 16'b0000010001100101;
            15'd12857: log10_cal = 16'b0000010001100101;
            15'd12858: log10_cal = 16'b0000010001100101;
            15'd12859: log10_cal = 16'b0000010001100101;
            15'd12860: log10_cal = 16'b0000010001100101;
            15'd12861: log10_cal = 16'b0000010001100101;
            15'd12862: log10_cal = 16'b0000010001100101;
            15'd12863: log10_cal = 16'b0000010001100101;
            15'd12864: log10_cal = 16'b0000010001100101;
            15'd12865: log10_cal = 16'b0000010001100101;
            15'd12866: log10_cal = 16'b0000010001100101;
            15'd12867: log10_cal = 16'b0000010001100101;
            15'd12868: log10_cal = 16'b0000010001100101;
            15'd12869: log10_cal = 16'b0000010001100101;
            15'd12870: log10_cal = 16'b0000010001100101;
            15'd12871: log10_cal = 16'b0000010001100101;
            15'd12872: log10_cal = 16'b0000010001100101;
            15'd12873: log10_cal = 16'b0000010001100101;
            15'd12874: log10_cal = 16'b0000010001100101;
            15'd12875: log10_cal = 16'b0000010001100101;
            15'd12876: log10_cal = 16'b0000010001100101;
            15'd12877: log10_cal = 16'b0000010001100101;
            15'd12878: log10_cal = 16'b0000010001100101;
            15'd12879: log10_cal = 16'b0000010001100101;
            15'd12880: log10_cal = 16'b0000010001100110;
            15'd12881: log10_cal = 16'b0000010001100110;
            15'd12882: log10_cal = 16'b0000010001100110;
            15'd12883: log10_cal = 16'b0000010001100110;
            15'd12884: log10_cal = 16'b0000010001100110;
            15'd12885: log10_cal = 16'b0000010001100110;
            15'd12886: log10_cal = 16'b0000010001100110;
            15'd12887: log10_cal = 16'b0000010001100110;
            15'd12888: log10_cal = 16'b0000010001100110;
            15'd12889: log10_cal = 16'b0000010001100110;
            15'd12890: log10_cal = 16'b0000010001100110;
            15'd12891: log10_cal = 16'b0000010001100110;
            15'd12892: log10_cal = 16'b0000010001100110;
            15'd12893: log10_cal = 16'b0000010001100110;
            15'd12894: log10_cal = 16'b0000010001100110;
            15'd12895: log10_cal = 16'b0000010001100110;
            15'd12896: log10_cal = 16'b0000010001100110;
            15'd12897: log10_cal = 16'b0000010001100110;
            15'd12898: log10_cal = 16'b0000010001100110;
            15'd12899: log10_cal = 16'b0000010001100110;
            15'd12900: log10_cal = 16'b0000010001100110;
            15'd12901: log10_cal = 16'b0000010001100110;
            15'd12902: log10_cal = 16'b0000010001100110;
            15'd12903: log10_cal = 16'b0000010001100110;
            15'd12904: log10_cal = 16'b0000010001100110;
            15'd12905: log10_cal = 16'b0000010001100110;
            15'd12906: log10_cal = 16'b0000010001100110;
            15'd12907: log10_cal = 16'b0000010001100110;
            15'd12908: log10_cal = 16'b0000010001100110;
            15'd12909: log10_cal = 16'b0000010001100111;
            15'd12910: log10_cal = 16'b0000010001100111;
            15'd12911: log10_cal = 16'b0000010001100111;
            15'd12912: log10_cal = 16'b0000010001100111;
            15'd12913: log10_cal = 16'b0000010001100111;
            15'd12914: log10_cal = 16'b0000010001100111;
            15'd12915: log10_cal = 16'b0000010001100111;
            15'd12916: log10_cal = 16'b0000010001100111;
            15'd12917: log10_cal = 16'b0000010001100111;
            15'd12918: log10_cal = 16'b0000010001100111;
            15'd12919: log10_cal = 16'b0000010001100111;
            15'd12920: log10_cal = 16'b0000010001100111;
            15'd12921: log10_cal = 16'b0000010001100111;
            15'd12922: log10_cal = 16'b0000010001100111;
            15'd12923: log10_cal = 16'b0000010001100111;
            15'd12924: log10_cal = 16'b0000010001100111;
            15'd12925: log10_cal = 16'b0000010001100111;
            15'd12926: log10_cal = 16'b0000010001100111;
            15'd12927: log10_cal = 16'b0000010001100111;
            15'd12928: log10_cal = 16'b0000010001100111;
            15'd12929: log10_cal = 16'b0000010001100111;
            15'd12930: log10_cal = 16'b0000010001100111;
            15'd12931: log10_cal = 16'b0000010001100111;
            15'd12932: log10_cal = 16'b0000010001100111;
            15'd12933: log10_cal = 16'b0000010001100111;
            15'd12934: log10_cal = 16'b0000010001100111;
            15'd12935: log10_cal = 16'b0000010001100111;
            15'd12936: log10_cal = 16'b0000010001100111;
            15'd12937: log10_cal = 16'b0000010001100111;
            15'd12938: log10_cal = 16'b0000010001101000;
            15'd12939: log10_cal = 16'b0000010001101000;
            15'd12940: log10_cal = 16'b0000010001101000;
            15'd12941: log10_cal = 16'b0000010001101000;
            15'd12942: log10_cal = 16'b0000010001101000;
            15'd12943: log10_cal = 16'b0000010001101000;
            15'd12944: log10_cal = 16'b0000010001101000;
            15'd12945: log10_cal = 16'b0000010001101000;
            15'd12946: log10_cal = 16'b0000010001101000;
            15'd12947: log10_cal = 16'b0000010001101000;
            15'd12948: log10_cal = 16'b0000010001101000;
            15'd12949: log10_cal = 16'b0000010001101000;
            15'd12950: log10_cal = 16'b0000010001101000;
            15'd12951: log10_cal = 16'b0000010001101000;
            15'd12952: log10_cal = 16'b0000010001101000;
            15'd12953: log10_cal = 16'b0000010001101000;
            15'd12954: log10_cal = 16'b0000010001101000;
            15'd12955: log10_cal = 16'b0000010001101000;
            15'd12956: log10_cal = 16'b0000010001101000;
            15'd12957: log10_cal = 16'b0000010001101000;
            15'd12958: log10_cal = 16'b0000010001101000;
            15'd12959: log10_cal = 16'b0000010001101000;
            15'd12960: log10_cal = 16'b0000010001101000;
            15'd12961: log10_cal = 16'b0000010001101000;
            15'd12962: log10_cal = 16'b0000010001101000;
            15'd12963: log10_cal = 16'b0000010001101000;
            15'd12964: log10_cal = 16'b0000010001101000;
            15'd12965: log10_cal = 16'b0000010001101000;
            15'd12966: log10_cal = 16'b0000010001101000;
            15'd12967: log10_cal = 16'b0000010001101001;
            15'd12968: log10_cal = 16'b0000010001101001;
            15'd12969: log10_cal = 16'b0000010001101001;
            15'd12970: log10_cal = 16'b0000010001101001;
            15'd12971: log10_cal = 16'b0000010001101001;
            15'd12972: log10_cal = 16'b0000010001101001;
            15'd12973: log10_cal = 16'b0000010001101001;
            15'd12974: log10_cal = 16'b0000010001101001;
            15'd12975: log10_cal = 16'b0000010001101001;
            15'd12976: log10_cal = 16'b0000010001101001;
            15'd12977: log10_cal = 16'b0000010001101001;
            15'd12978: log10_cal = 16'b0000010001101001;
            15'd12979: log10_cal = 16'b0000010001101001;
            15'd12980: log10_cal = 16'b0000010001101001;
            15'd12981: log10_cal = 16'b0000010001101001;
            15'd12982: log10_cal = 16'b0000010001101001;
            15'd12983: log10_cal = 16'b0000010001101001;
            15'd12984: log10_cal = 16'b0000010001101001;
            15'd12985: log10_cal = 16'b0000010001101001;
            15'd12986: log10_cal = 16'b0000010001101001;
            15'd12987: log10_cal = 16'b0000010001101001;
            15'd12988: log10_cal = 16'b0000010001101001;
            15'd12989: log10_cal = 16'b0000010001101001;
            15'd12990: log10_cal = 16'b0000010001101001;
            15'd12991: log10_cal = 16'b0000010001101001;
            15'd12992: log10_cal = 16'b0000010001101001;
            15'd12993: log10_cal = 16'b0000010001101001;
            15'd12994: log10_cal = 16'b0000010001101001;
            15'd12995: log10_cal = 16'b0000010001101001;
            15'd12996: log10_cal = 16'b0000010001101001;
            15'd12997: log10_cal = 16'b0000010001101010;
            15'd12998: log10_cal = 16'b0000010001101010;
            15'd12999: log10_cal = 16'b0000010001101010;
            15'd13000: log10_cal = 16'b0000010001101010;
            15'd13001: log10_cal = 16'b0000010001101010;
            15'd13002: log10_cal = 16'b0000010001101010;
            15'd13003: log10_cal = 16'b0000010001101010;
            15'd13004: log10_cal = 16'b0000010001101010;
            15'd13005: log10_cal = 16'b0000010001101010;
            15'd13006: log10_cal = 16'b0000010001101010;
            15'd13007: log10_cal = 16'b0000010001101010;
            15'd13008: log10_cal = 16'b0000010001101010;
            15'd13009: log10_cal = 16'b0000010001101010;
            15'd13010: log10_cal = 16'b0000010001101010;
            15'd13011: log10_cal = 16'b0000010001101010;
            15'd13012: log10_cal = 16'b0000010001101010;
            15'd13013: log10_cal = 16'b0000010001101010;
            15'd13014: log10_cal = 16'b0000010001101010;
            15'd13015: log10_cal = 16'b0000010001101010;
            15'd13016: log10_cal = 16'b0000010001101010;
            15'd13017: log10_cal = 16'b0000010001101010;
            15'd13018: log10_cal = 16'b0000010001101010;
            15'd13019: log10_cal = 16'b0000010001101010;
            15'd13020: log10_cal = 16'b0000010001101010;
            15'd13021: log10_cal = 16'b0000010001101010;
            15'd13022: log10_cal = 16'b0000010001101010;
            15'd13023: log10_cal = 16'b0000010001101010;
            15'd13024: log10_cal = 16'b0000010001101010;
            15'd13025: log10_cal = 16'b0000010001101010;
            15'd13026: log10_cal = 16'b0000010001101011;
            15'd13027: log10_cal = 16'b0000010001101011;
            15'd13028: log10_cal = 16'b0000010001101011;
            15'd13029: log10_cal = 16'b0000010001101011;
            15'd13030: log10_cal = 16'b0000010001101011;
            15'd13031: log10_cal = 16'b0000010001101011;
            15'd13032: log10_cal = 16'b0000010001101011;
            15'd13033: log10_cal = 16'b0000010001101011;
            15'd13034: log10_cal = 16'b0000010001101011;
            15'd13035: log10_cal = 16'b0000010001101011;
            15'd13036: log10_cal = 16'b0000010001101011;
            15'd13037: log10_cal = 16'b0000010001101011;
            15'd13038: log10_cal = 16'b0000010001101011;
            15'd13039: log10_cal = 16'b0000010001101011;
            15'd13040: log10_cal = 16'b0000010001101011;
            15'd13041: log10_cal = 16'b0000010001101011;
            15'd13042: log10_cal = 16'b0000010001101011;
            15'd13043: log10_cal = 16'b0000010001101011;
            15'd13044: log10_cal = 16'b0000010001101011;
            15'd13045: log10_cal = 16'b0000010001101011;
            15'd13046: log10_cal = 16'b0000010001101011;
            15'd13047: log10_cal = 16'b0000010001101011;
            15'd13048: log10_cal = 16'b0000010001101011;
            15'd13049: log10_cal = 16'b0000010001101011;
            15'd13050: log10_cal = 16'b0000010001101011;
            15'd13051: log10_cal = 16'b0000010001101011;
            15'd13052: log10_cal = 16'b0000010001101011;
            15'd13053: log10_cal = 16'b0000010001101011;
            15'd13054: log10_cal = 16'b0000010001101011;
            15'd13055: log10_cal = 16'b0000010001101100;
            15'd13056: log10_cal = 16'b0000010001101100;
            15'd13057: log10_cal = 16'b0000010001101100;
            15'd13058: log10_cal = 16'b0000010001101100;
            15'd13059: log10_cal = 16'b0000010001101100;
            15'd13060: log10_cal = 16'b0000010001101100;
            15'd13061: log10_cal = 16'b0000010001101100;
            15'd13062: log10_cal = 16'b0000010001101100;
            15'd13063: log10_cal = 16'b0000010001101100;
            15'd13064: log10_cal = 16'b0000010001101100;
            15'd13065: log10_cal = 16'b0000010001101100;
            15'd13066: log10_cal = 16'b0000010001101100;
            15'd13067: log10_cal = 16'b0000010001101100;
            15'd13068: log10_cal = 16'b0000010001101100;
            15'd13069: log10_cal = 16'b0000010001101100;
            15'd13070: log10_cal = 16'b0000010001101100;
            15'd13071: log10_cal = 16'b0000010001101100;
            15'd13072: log10_cal = 16'b0000010001101100;
            15'd13073: log10_cal = 16'b0000010001101100;
            15'd13074: log10_cal = 16'b0000010001101100;
            15'd13075: log10_cal = 16'b0000010001101100;
            15'd13076: log10_cal = 16'b0000010001101100;
            15'd13077: log10_cal = 16'b0000010001101100;
            15'd13078: log10_cal = 16'b0000010001101100;
            15'd13079: log10_cal = 16'b0000010001101100;
            15'd13080: log10_cal = 16'b0000010001101100;
            15'd13081: log10_cal = 16'b0000010001101100;
            15'd13082: log10_cal = 16'b0000010001101100;
            15'd13083: log10_cal = 16'b0000010001101100;
            15'd13084: log10_cal = 16'b0000010001101100;
            15'd13085: log10_cal = 16'b0000010001101101;
            15'd13086: log10_cal = 16'b0000010001101101;
            15'd13087: log10_cal = 16'b0000010001101101;
            15'd13088: log10_cal = 16'b0000010001101101;
            15'd13089: log10_cal = 16'b0000010001101101;
            15'd13090: log10_cal = 16'b0000010001101101;
            15'd13091: log10_cal = 16'b0000010001101101;
            15'd13092: log10_cal = 16'b0000010001101101;
            15'd13093: log10_cal = 16'b0000010001101101;
            15'd13094: log10_cal = 16'b0000010001101101;
            15'd13095: log10_cal = 16'b0000010001101101;
            15'd13096: log10_cal = 16'b0000010001101101;
            15'd13097: log10_cal = 16'b0000010001101101;
            15'd13098: log10_cal = 16'b0000010001101101;
            15'd13099: log10_cal = 16'b0000010001101101;
            15'd13100: log10_cal = 16'b0000010001101101;
            15'd13101: log10_cal = 16'b0000010001101101;
            15'd13102: log10_cal = 16'b0000010001101101;
            15'd13103: log10_cal = 16'b0000010001101101;
            15'd13104: log10_cal = 16'b0000010001101101;
            15'd13105: log10_cal = 16'b0000010001101101;
            15'd13106: log10_cal = 16'b0000010001101101;
            15'd13107: log10_cal = 16'b0000010001101101;
            15'd13108: log10_cal = 16'b0000010001101101;
            15'd13109: log10_cal = 16'b0000010001101101;
            15'd13110: log10_cal = 16'b0000010001101101;
            15'd13111: log10_cal = 16'b0000010001101101;
            15'd13112: log10_cal = 16'b0000010001101101;
            15'd13113: log10_cal = 16'b0000010001101101;
            15'd13114: log10_cal = 16'b0000010001101110;
            15'd13115: log10_cal = 16'b0000010001101110;
            15'd13116: log10_cal = 16'b0000010001101110;
            15'd13117: log10_cal = 16'b0000010001101110;
            15'd13118: log10_cal = 16'b0000010001101110;
            15'd13119: log10_cal = 16'b0000010001101110;
            15'd13120: log10_cal = 16'b0000010001101110;
            15'd13121: log10_cal = 16'b0000010001101110;
            15'd13122: log10_cal = 16'b0000010001101110;
            15'd13123: log10_cal = 16'b0000010001101110;
            15'd13124: log10_cal = 16'b0000010001101110;
            15'd13125: log10_cal = 16'b0000010001101110;
            15'd13126: log10_cal = 16'b0000010001101110;
            15'd13127: log10_cal = 16'b0000010001101110;
            15'd13128: log10_cal = 16'b0000010001101110;
            15'd13129: log10_cal = 16'b0000010001101110;
            15'd13130: log10_cal = 16'b0000010001101110;
            15'd13131: log10_cal = 16'b0000010001101110;
            15'd13132: log10_cal = 16'b0000010001101110;
            15'd13133: log10_cal = 16'b0000010001101110;
            15'd13134: log10_cal = 16'b0000010001101110;
            15'd13135: log10_cal = 16'b0000010001101110;
            15'd13136: log10_cal = 16'b0000010001101110;
            15'd13137: log10_cal = 16'b0000010001101110;
            15'd13138: log10_cal = 16'b0000010001101110;
            15'd13139: log10_cal = 16'b0000010001101110;
            15'd13140: log10_cal = 16'b0000010001101110;
            15'd13141: log10_cal = 16'b0000010001101110;
            15'd13142: log10_cal = 16'b0000010001101110;
            15'd13143: log10_cal = 16'b0000010001101110;
            15'd13144: log10_cal = 16'b0000010001101111;
            15'd13145: log10_cal = 16'b0000010001101111;
            15'd13146: log10_cal = 16'b0000010001101111;
            15'd13147: log10_cal = 16'b0000010001101111;
            15'd13148: log10_cal = 16'b0000010001101111;
            15'd13149: log10_cal = 16'b0000010001101111;
            15'd13150: log10_cal = 16'b0000010001101111;
            15'd13151: log10_cal = 16'b0000010001101111;
            15'd13152: log10_cal = 16'b0000010001101111;
            15'd13153: log10_cal = 16'b0000010001101111;
            15'd13154: log10_cal = 16'b0000010001101111;
            15'd13155: log10_cal = 16'b0000010001101111;
            15'd13156: log10_cal = 16'b0000010001101111;
            15'd13157: log10_cal = 16'b0000010001101111;
            15'd13158: log10_cal = 16'b0000010001101111;
            15'd13159: log10_cal = 16'b0000010001101111;
            15'd13160: log10_cal = 16'b0000010001101111;
            15'd13161: log10_cal = 16'b0000010001101111;
            15'd13162: log10_cal = 16'b0000010001101111;
            15'd13163: log10_cal = 16'b0000010001101111;
            15'd13164: log10_cal = 16'b0000010001101111;
            15'd13165: log10_cal = 16'b0000010001101111;
            15'd13166: log10_cal = 16'b0000010001101111;
            15'd13167: log10_cal = 16'b0000010001101111;
            15'd13168: log10_cal = 16'b0000010001101111;
            15'd13169: log10_cal = 16'b0000010001101111;
            15'd13170: log10_cal = 16'b0000010001101111;
            15'd13171: log10_cal = 16'b0000010001101111;
            15'd13172: log10_cal = 16'b0000010001101111;
            15'd13173: log10_cal = 16'b0000010001110000;
            15'd13174: log10_cal = 16'b0000010001110000;
            15'd13175: log10_cal = 16'b0000010001110000;
            15'd13176: log10_cal = 16'b0000010001110000;
            15'd13177: log10_cal = 16'b0000010001110000;
            15'd13178: log10_cal = 16'b0000010001110000;
            15'd13179: log10_cal = 16'b0000010001110000;
            15'd13180: log10_cal = 16'b0000010001110000;
            15'd13181: log10_cal = 16'b0000010001110000;
            15'd13182: log10_cal = 16'b0000010001110000;
            15'd13183: log10_cal = 16'b0000010001110000;
            15'd13184: log10_cal = 16'b0000010001110000;
            15'd13185: log10_cal = 16'b0000010001110000;
            15'd13186: log10_cal = 16'b0000010001110000;
            15'd13187: log10_cal = 16'b0000010001110000;
            15'd13188: log10_cal = 16'b0000010001110000;
            15'd13189: log10_cal = 16'b0000010001110000;
            15'd13190: log10_cal = 16'b0000010001110000;
            15'd13191: log10_cal = 16'b0000010001110000;
            15'd13192: log10_cal = 16'b0000010001110000;
            15'd13193: log10_cal = 16'b0000010001110000;
            15'd13194: log10_cal = 16'b0000010001110000;
            15'd13195: log10_cal = 16'b0000010001110000;
            15'd13196: log10_cal = 16'b0000010001110000;
            15'd13197: log10_cal = 16'b0000010001110000;
            15'd13198: log10_cal = 16'b0000010001110000;
            15'd13199: log10_cal = 16'b0000010001110000;
            15'd13200: log10_cal = 16'b0000010001110000;
            15'd13201: log10_cal = 16'b0000010001110000;
            15'd13202: log10_cal = 16'b0000010001110000;
            15'd13203: log10_cal = 16'b0000010001110001;
            15'd13204: log10_cal = 16'b0000010001110001;
            15'd13205: log10_cal = 16'b0000010001110001;
            15'd13206: log10_cal = 16'b0000010001110001;
            15'd13207: log10_cal = 16'b0000010001110001;
            15'd13208: log10_cal = 16'b0000010001110001;
            15'd13209: log10_cal = 16'b0000010001110001;
            15'd13210: log10_cal = 16'b0000010001110001;
            15'd13211: log10_cal = 16'b0000010001110001;
            15'd13212: log10_cal = 16'b0000010001110001;
            15'd13213: log10_cal = 16'b0000010001110001;
            15'd13214: log10_cal = 16'b0000010001110001;
            15'd13215: log10_cal = 16'b0000010001110001;
            15'd13216: log10_cal = 16'b0000010001110001;
            15'd13217: log10_cal = 16'b0000010001110001;
            15'd13218: log10_cal = 16'b0000010001110001;
            15'd13219: log10_cal = 16'b0000010001110001;
            15'd13220: log10_cal = 16'b0000010001110001;
            15'd13221: log10_cal = 16'b0000010001110001;
            15'd13222: log10_cal = 16'b0000010001110001;
            15'd13223: log10_cal = 16'b0000010001110001;
            15'd13224: log10_cal = 16'b0000010001110001;
            15'd13225: log10_cal = 16'b0000010001110001;
            15'd13226: log10_cal = 16'b0000010001110001;
            15'd13227: log10_cal = 16'b0000010001110001;
            15'd13228: log10_cal = 16'b0000010001110001;
            15'd13229: log10_cal = 16'b0000010001110001;
            15'd13230: log10_cal = 16'b0000010001110001;
            15'd13231: log10_cal = 16'b0000010001110001;
            15'd13232: log10_cal = 16'b0000010001110001;
            15'd13233: log10_cal = 16'b0000010001110010;
            15'd13234: log10_cal = 16'b0000010001110010;
            15'd13235: log10_cal = 16'b0000010001110010;
            15'd13236: log10_cal = 16'b0000010001110010;
            15'd13237: log10_cal = 16'b0000010001110010;
            15'd13238: log10_cal = 16'b0000010001110010;
            15'd13239: log10_cal = 16'b0000010001110010;
            15'd13240: log10_cal = 16'b0000010001110010;
            15'd13241: log10_cal = 16'b0000010001110010;
            15'd13242: log10_cal = 16'b0000010001110010;
            15'd13243: log10_cal = 16'b0000010001110010;
            15'd13244: log10_cal = 16'b0000010001110010;
            15'd13245: log10_cal = 16'b0000010001110010;
            15'd13246: log10_cal = 16'b0000010001110010;
            15'd13247: log10_cal = 16'b0000010001110010;
            15'd13248: log10_cal = 16'b0000010001110010;
            15'd13249: log10_cal = 16'b0000010001110010;
            15'd13250: log10_cal = 16'b0000010001110010;
            15'd13251: log10_cal = 16'b0000010001110010;
            15'd13252: log10_cal = 16'b0000010001110010;
            15'd13253: log10_cal = 16'b0000010001110010;
            15'd13254: log10_cal = 16'b0000010001110010;
            15'd13255: log10_cal = 16'b0000010001110010;
            15'd13256: log10_cal = 16'b0000010001110010;
            15'd13257: log10_cal = 16'b0000010001110010;
            15'd13258: log10_cal = 16'b0000010001110010;
            15'd13259: log10_cal = 16'b0000010001110010;
            15'd13260: log10_cal = 16'b0000010001110010;
            15'd13261: log10_cal = 16'b0000010001110010;
            15'd13262: log10_cal = 16'b0000010001110011;
            15'd13263: log10_cal = 16'b0000010001110011;
            15'd13264: log10_cal = 16'b0000010001110011;
            15'd13265: log10_cal = 16'b0000010001110011;
            15'd13266: log10_cal = 16'b0000010001110011;
            15'd13267: log10_cal = 16'b0000010001110011;
            15'd13268: log10_cal = 16'b0000010001110011;
            15'd13269: log10_cal = 16'b0000010001110011;
            15'd13270: log10_cal = 16'b0000010001110011;
            15'd13271: log10_cal = 16'b0000010001110011;
            15'd13272: log10_cal = 16'b0000010001110011;
            15'd13273: log10_cal = 16'b0000010001110011;
            15'd13274: log10_cal = 16'b0000010001110011;
            15'd13275: log10_cal = 16'b0000010001110011;
            15'd13276: log10_cal = 16'b0000010001110011;
            15'd13277: log10_cal = 16'b0000010001110011;
            15'd13278: log10_cal = 16'b0000010001110011;
            15'd13279: log10_cal = 16'b0000010001110011;
            15'd13280: log10_cal = 16'b0000010001110011;
            15'd13281: log10_cal = 16'b0000010001110011;
            15'd13282: log10_cal = 16'b0000010001110011;
            15'd13283: log10_cal = 16'b0000010001110011;
            15'd13284: log10_cal = 16'b0000010001110011;
            15'd13285: log10_cal = 16'b0000010001110011;
            15'd13286: log10_cal = 16'b0000010001110011;
            15'd13287: log10_cal = 16'b0000010001110011;
            15'd13288: log10_cal = 16'b0000010001110011;
            15'd13289: log10_cal = 16'b0000010001110011;
            15'd13290: log10_cal = 16'b0000010001110011;
            15'd13291: log10_cal = 16'b0000010001110011;
            15'd13292: log10_cal = 16'b0000010001110100;
            15'd13293: log10_cal = 16'b0000010001110100;
            15'd13294: log10_cal = 16'b0000010001110100;
            15'd13295: log10_cal = 16'b0000010001110100;
            15'd13296: log10_cal = 16'b0000010001110100;
            15'd13297: log10_cal = 16'b0000010001110100;
            15'd13298: log10_cal = 16'b0000010001110100;
            15'd13299: log10_cal = 16'b0000010001110100;
            15'd13300: log10_cal = 16'b0000010001110100;
            15'd13301: log10_cal = 16'b0000010001110100;
            15'd13302: log10_cal = 16'b0000010001110100;
            15'd13303: log10_cal = 16'b0000010001110100;
            15'd13304: log10_cal = 16'b0000010001110100;
            15'd13305: log10_cal = 16'b0000010001110100;
            15'd13306: log10_cal = 16'b0000010001110100;
            15'd13307: log10_cal = 16'b0000010001110100;
            15'd13308: log10_cal = 16'b0000010001110100;
            15'd13309: log10_cal = 16'b0000010001110100;
            15'd13310: log10_cal = 16'b0000010001110100;
            15'd13311: log10_cal = 16'b0000010001110100;
            15'd13312: log10_cal = 16'b0000010001110100;
            15'd13313: log10_cal = 16'b0000010001110100;
            15'd13314: log10_cal = 16'b0000010001110100;
            15'd13315: log10_cal = 16'b0000010001110100;
            15'd13316: log10_cal = 16'b0000010001110100;
            15'd13317: log10_cal = 16'b0000010001110100;
            15'd13318: log10_cal = 16'b0000010001110100;
            15'd13319: log10_cal = 16'b0000010001110100;
            15'd13320: log10_cal = 16'b0000010001110100;
            15'd13321: log10_cal = 16'b0000010001110100;
            15'd13322: log10_cal = 16'b0000010001110101;
            15'd13323: log10_cal = 16'b0000010001110101;
            15'd13324: log10_cal = 16'b0000010001110101;
            15'd13325: log10_cal = 16'b0000010001110101;
            15'd13326: log10_cal = 16'b0000010001110101;
            15'd13327: log10_cal = 16'b0000010001110101;
            15'd13328: log10_cal = 16'b0000010001110101;
            15'd13329: log10_cal = 16'b0000010001110101;
            15'd13330: log10_cal = 16'b0000010001110101;
            15'd13331: log10_cal = 16'b0000010001110101;
            15'd13332: log10_cal = 16'b0000010001110101;
            15'd13333: log10_cal = 16'b0000010001110101;
            15'd13334: log10_cal = 16'b0000010001110101;
            15'd13335: log10_cal = 16'b0000010001110101;
            15'd13336: log10_cal = 16'b0000010001110101;
            15'd13337: log10_cal = 16'b0000010001110101;
            15'd13338: log10_cal = 16'b0000010001110101;
            15'd13339: log10_cal = 16'b0000010001110101;
            15'd13340: log10_cal = 16'b0000010001110101;
            15'd13341: log10_cal = 16'b0000010001110101;
            15'd13342: log10_cal = 16'b0000010001110101;
            15'd13343: log10_cal = 16'b0000010001110101;
            15'd13344: log10_cal = 16'b0000010001110101;
            15'd13345: log10_cal = 16'b0000010001110101;
            15'd13346: log10_cal = 16'b0000010001110101;
            15'd13347: log10_cal = 16'b0000010001110101;
            15'd13348: log10_cal = 16'b0000010001110101;
            15'd13349: log10_cal = 16'b0000010001110101;
            15'd13350: log10_cal = 16'b0000010001110101;
            15'd13351: log10_cal = 16'b0000010001110101;
            15'd13352: log10_cal = 16'b0000010001110110;
            15'd13353: log10_cal = 16'b0000010001110110;
            15'd13354: log10_cal = 16'b0000010001110110;
            15'd13355: log10_cal = 16'b0000010001110110;
            15'd13356: log10_cal = 16'b0000010001110110;
            15'd13357: log10_cal = 16'b0000010001110110;
            15'd13358: log10_cal = 16'b0000010001110110;
            15'd13359: log10_cal = 16'b0000010001110110;
            15'd13360: log10_cal = 16'b0000010001110110;
            15'd13361: log10_cal = 16'b0000010001110110;
            15'd13362: log10_cal = 16'b0000010001110110;
            15'd13363: log10_cal = 16'b0000010001110110;
            15'd13364: log10_cal = 16'b0000010001110110;
            15'd13365: log10_cal = 16'b0000010001110110;
            15'd13366: log10_cal = 16'b0000010001110110;
            15'd13367: log10_cal = 16'b0000010001110110;
            15'd13368: log10_cal = 16'b0000010001110110;
            15'd13369: log10_cal = 16'b0000010001110110;
            15'd13370: log10_cal = 16'b0000010001110110;
            15'd13371: log10_cal = 16'b0000010001110110;
            15'd13372: log10_cal = 16'b0000010001110110;
            15'd13373: log10_cal = 16'b0000010001110110;
            15'd13374: log10_cal = 16'b0000010001110110;
            15'd13375: log10_cal = 16'b0000010001110110;
            15'd13376: log10_cal = 16'b0000010001110110;
            15'd13377: log10_cal = 16'b0000010001110110;
            15'd13378: log10_cal = 16'b0000010001110110;
            15'd13379: log10_cal = 16'b0000010001110110;
            15'd13380: log10_cal = 16'b0000010001110110;
            15'd13381: log10_cal = 16'b0000010001110110;
            15'd13382: log10_cal = 16'b0000010001110111;
            15'd13383: log10_cal = 16'b0000010001110111;
            15'd13384: log10_cal = 16'b0000010001110111;
            15'd13385: log10_cal = 16'b0000010001110111;
            15'd13386: log10_cal = 16'b0000010001110111;
            15'd13387: log10_cal = 16'b0000010001110111;
            15'd13388: log10_cal = 16'b0000010001110111;
            15'd13389: log10_cal = 16'b0000010001110111;
            15'd13390: log10_cal = 16'b0000010001110111;
            15'd13391: log10_cal = 16'b0000010001110111;
            15'd13392: log10_cal = 16'b0000010001110111;
            15'd13393: log10_cal = 16'b0000010001110111;
            15'd13394: log10_cal = 16'b0000010001110111;
            15'd13395: log10_cal = 16'b0000010001110111;
            15'd13396: log10_cal = 16'b0000010001110111;
            15'd13397: log10_cal = 16'b0000010001110111;
            15'd13398: log10_cal = 16'b0000010001110111;
            15'd13399: log10_cal = 16'b0000010001110111;
            15'd13400: log10_cal = 16'b0000010001110111;
            15'd13401: log10_cal = 16'b0000010001110111;
            15'd13402: log10_cal = 16'b0000010001110111;
            15'd13403: log10_cal = 16'b0000010001110111;
            15'd13404: log10_cal = 16'b0000010001110111;
            15'd13405: log10_cal = 16'b0000010001110111;
            15'd13406: log10_cal = 16'b0000010001110111;
            15'd13407: log10_cal = 16'b0000010001110111;
            15'd13408: log10_cal = 16'b0000010001110111;
            15'd13409: log10_cal = 16'b0000010001110111;
            15'd13410: log10_cal = 16'b0000010001110111;
            15'd13411: log10_cal = 16'b0000010001110111;
            15'd13412: log10_cal = 16'b0000010001111000;
            15'd13413: log10_cal = 16'b0000010001111000;
            15'd13414: log10_cal = 16'b0000010001111000;
            15'd13415: log10_cal = 16'b0000010001111000;
            15'd13416: log10_cal = 16'b0000010001111000;
            15'd13417: log10_cal = 16'b0000010001111000;
            15'd13418: log10_cal = 16'b0000010001111000;
            15'd13419: log10_cal = 16'b0000010001111000;
            15'd13420: log10_cal = 16'b0000010001111000;
            15'd13421: log10_cal = 16'b0000010001111000;
            15'd13422: log10_cal = 16'b0000010001111000;
            15'd13423: log10_cal = 16'b0000010001111000;
            15'd13424: log10_cal = 16'b0000010001111000;
            15'd13425: log10_cal = 16'b0000010001111000;
            15'd13426: log10_cal = 16'b0000010001111000;
            15'd13427: log10_cal = 16'b0000010001111000;
            15'd13428: log10_cal = 16'b0000010001111000;
            15'd13429: log10_cal = 16'b0000010001111000;
            15'd13430: log10_cal = 16'b0000010001111000;
            15'd13431: log10_cal = 16'b0000010001111000;
            15'd13432: log10_cal = 16'b0000010001111000;
            15'd13433: log10_cal = 16'b0000010001111000;
            15'd13434: log10_cal = 16'b0000010001111000;
            15'd13435: log10_cal = 16'b0000010001111000;
            15'd13436: log10_cal = 16'b0000010001111000;
            15'd13437: log10_cal = 16'b0000010001111000;
            15'd13438: log10_cal = 16'b0000010001111000;
            15'd13439: log10_cal = 16'b0000010001111000;
            15'd13440: log10_cal = 16'b0000010001111000;
            15'd13441: log10_cal = 16'b0000010001111000;
            15'd13442: log10_cal = 16'b0000010001111000;
            15'd13443: log10_cal = 16'b0000010001111001;
            15'd13444: log10_cal = 16'b0000010001111001;
            15'd13445: log10_cal = 16'b0000010001111001;
            15'd13446: log10_cal = 16'b0000010001111001;
            15'd13447: log10_cal = 16'b0000010001111001;
            15'd13448: log10_cal = 16'b0000010001111001;
            15'd13449: log10_cal = 16'b0000010001111001;
            15'd13450: log10_cal = 16'b0000010001111001;
            15'd13451: log10_cal = 16'b0000010001111001;
            15'd13452: log10_cal = 16'b0000010001111001;
            15'd13453: log10_cal = 16'b0000010001111001;
            15'd13454: log10_cal = 16'b0000010001111001;
            15'd13455: log10_cal = 16'b0000010001111001;
            15'd13456: log10_cal = 16'b0000010001111001;
            15'd13457: log10_cal = 16'b0000010001111001;
            15'd13458: log10_cal = 16'b0000010001111001;
            15'd13459: log10_cal = 16'b0000010001111001;
            15'd13460: log10_cal = 16'b0000010001111001;
            15'd13461: log10_cal = 16'b0000010001111001;
            15'd13462: log10_cal = 16'b0000010001111001;
            15'd13463: log10_cal = 16'b0000010001111001;
            15'd13464: log10_cal = 16'b0000010001111001;
            15'd13465: log10_cal = 16'b0000010001111001;
            15'd13466: log10_cal = 16'b0000010001111001;
            15'd13467: log10_cal = 16'b0000010001111001;
            15'd13468: log10_cal = 16'b0000010001111001;
            15'd13469: log10_cal = 16'b0000010001111001;
            15'd13470: log10_cal = 16'b0000010001111001;
            15'd13471: log10_cal = 16'b0000010001111001;
            15'd13472: log10_cal = 16'b0000010001111001;
            15'd13473: log10_cal = 16'b0000010001111010;
            15'd13474: log10_cal = 16'b0000010001111010;
            15'd13475: log10_cal = 16'b0000010001111010;
            15'd13476: log10_cal = 16'b0000010001111010;
            15'd13477: log10_cal = 16'b0000010001111010;
            15'd13478: log10_cal = 16'b0000010001111010;
            15'd13479: log10_cal = 16'b0000010001111010;
            15'd13480: log10_cal = 16'b0000010001111010;
            15'd13481: log10_cal = 16'b0000010001111010;
            15'd13482: log10_cal = 16'b0000010001111010;
            15'd13483: log10_cal = 16'b0000010001111010;
            15'd13484: log10_cal = 16'b0000010001111010;
            15'd13485: log10_cal = 16'b0000010001111010;
            15'd13486: log10_cal = 16'b0000010001111010;
            15'd13487: log10_cal = 16'b0000010001111010;
            15'd13488: log10_cal = 16'b0000010001111010;
            15'd13489: log10_cal = 16'b0000010001111010;
            15'd13490: log10_cal = 16'b0000010001111010;
            15'd13491: log10_cal = 16'b0000010001111010;
            15'd13492: log10_cal = 16'b0000010001111010;
            15'd13493: log10_cal = 16'b0000010001111010;
            15'd13494: log10_cal = 16'b0000010001111010;
            15'd13495: log10_cal = 16'b0000010001111010;
            15'd13496: log10_cal = 16'b0000010001111010;
            15'd13497: log10_cal = 16'b0000010001111010;
            15'd13498: log10_cal = 16'b0000010001111010;
            15'd13499: log10_cal = 16'b0000010001111010;
            15'd13500: log10_cal = 16'b0000010001111010;
            15'd13501: log10_cal = 16'b0000010001111010;
            15'd13502: log10_cal = 16'b0000010001111010;
            15'd13503: log10_cal = 16'b0000010001111011;
            15'd13504: log10_cal = 16'b0000010001111011;
            15'd13505: log10_cal = 16'b0000010001111011;
            15'd13506: log10_cal = 16'b0000010001111011;
            15'd13507: log10_cal = 16'b0000010001111011;
            15'd13508: log10_cal = 16'b0000010001111011;
            15'd13509: log10_cal = 16'b0000010001111011;
            15'd13510: log10_cal = 16'b0000010001111011;
            15'd13511: log10_cal = 16'b0000010001111011;
            15'd13512: log10_cal = 16'b0000010001111011;
            15'd13513: log10_cal = 16'b0000010001111011;
            15'd13514: log10_cal = 16'b0000010001111011;
            15'd13515: log10_cal = 16'b0000010001111011;
            15'd13516: log10_cal = 16'b0000010001111011;
            15'd13517: log10_cal = 16'b0000010001111011;
            15'd13518: log10_cal = 16'b0000010001111011;
            15'd13519: log10_cal = 16'b0000010001111011;
            15'd13520: log10_cal = 16'b0000010001111011;
            15'd13521: log10_cal = 16'b0000010001111011;
            15'd13522: log10_cal = 16'b0000010001111011;
            15'd13523: log10_cal = 16'b0000010001111011;
            15'd13524: log10_cal = 16'b0000010001111011;
            15'd13525: log10_cal = 16'b0000010001111011;
            15'd13526: log10_cal = 16'b0000010001111011;
            15'd13527: log10_cal = 16'b0000010001111011;
            15'd13528: log10_cal = 16'b0000010001111011;
            15'd13529: log10_cal = 16'b0000010001111011;
            15'd13530: log10_cal = 16'b0000010001111011;
            15'd13531: log10_cal = 16'b0000010001111011;
            15'd13532: log10_cal = 16'b0000010001111011;
            15'd13533: log10_cal = 16'b0000010001111100;
            15'd13534: log10_cal = 16'b0000010001111100;
            15'd13535: log10_cal = 16'b0000010001111100;
            15'd13536: log10_cal = 16'b0000010001111100;
            15'd13537: log10_cal = 16'b0000010001111100;
            15'd13538: log10_cal = 16'b0000010001111100;
            15'd13539: log10_cal = 16'b0000010001111100;
            15'd13540: log10_cal = 16'b0000010001111100;
            15'd13541: log10_cal = 16'b0000010001111100;
            15'd13542: log10_cal = 16'b0000010001111100;
            15'd13543: log10_cal = 16'b0000010001111100;
            15'd13544: log10_cal = 16'b0000010001111100;
            15'd13545: log10_cal = 16'b0000010001111100;
            15'd13546: log10_cal = 16'b0000010001111100;
            15'd13547: log10_cal = 16'b0000010001111100;
            15'd13548: log10_cal = 16'b0000010001111100;
            15'd13549: log10_cal = 16'b0000010001111100;
            15'd13550: log10_cal = 16'b0000010001111100;
            15'd13551: log10_cal = 16'b0000010001111100;
            15'd13552: log10_cal = 16'b0000010001111100;
            15'd13553: log10_cal = 16'b0000010001111100;
            15'd13554: log10_cal = 16'b0000010001111100;
            15'd13555: log10_cal = 16'b0000010001111100;
            15'd13556: log10_cal = 16'b0000010001111100;
            15'd13557: log10_cal = 16'b0000010001111100;
            15'd13558: log10_cal = 16'b0000010001111100;
            15'd13559: log10_cal = 16'b0000010001111100;
            15'd13560: log10_cal = 16'b0000010001111100;
            15'd13561: log10_cal = 16'b0000010001111100;
            15'd13562: log10_cal = 16'b0000010001111100;
            15'd13563: log10_cal = 16'b0000010001111100;
            15'd13564: log10_cal = 16'b0000010001111101;
            15'd13565: log10_cal = 16'b0000010001111101;
            15'd13566: log10_cal = 16'b0000010001111101;
            15'd13567: log10_cal = 16'b0000010001111101;
            15'd13568: log10_cal = 16'b0000010001111101;
            15'd13569: log10_cal = 16'b0000010001111101;
            15'd13570: log10_cal = 16'b0000010001111101;
            15'd13571: log10_cal = 16'b0000010001111101;
            15'd13572: log10_cal = 16'b0000010001111101;
            15'd13573: log10_cal = 16'b0000010001111101;
            15'd13574: log10_cal = 16'b0000010001111101;
            15'd13575: log10_cal = 16'b0000010001111101;
            15'd13576: log10_cal = 16'b0000010001111101;
            15'd13577: log10_cal = 16'b0000010001111101;
            15'd13578: log10_cal = 16'b0000010001111101;
            15'd13579: log10_cal = 16'b0000010001111101;
            15'd13580: log10_cal = 16'b0000010001111101;
            15'd13581: log10_cal = 16'b0000010001111101;
            15'd13582: log10_cal = 16'b0000010001111101;
            15'd13583: log10_cal = 16'b0000010001111101;
            15'd13584: log10_cal = 16'b0000010001111101;
            15'd13585: log10_cal = 16'b0000010001111101;
            15'd13586: log10_cal = 16'b0000010001111101;
            15'd13587: log10_cal = 16'b0000010001111101;
            15'd13588: log10_cal = 16'b0000010001111101;
            15'd13589: log10_cal = 16'b0000010001111101;
            15'd13590: log10_cal = 16'b0000010001111101;
            15'd13591: log10_cal = 16'b0000010001111101;
            15'd13592: log10_cal = 16'b0000010001111101;
            15'd13593: log10_cal = 16'b0000010001111101;
            15'd13594: log10_cal = 16'b0000010001111110;
            15'd13595: log10_cal = 16'b0000010001111110;
            15'd13596: log10_cal = 16'b0000010001111110;
            15'd13597: log10_cal = 16'b0000010001111110;
            15'd13598: log10_cal = 16'b0000010001111110;
            15'd13599: log10_cal = 16'b0000010001111110;
            15'd13600: log10_cal = 16'b0000010001111110;
            15'd13601: log10_cal = 16'b0000010001111110;
            15'd13602: log10_cal = 16'b0000010001111110;
            15'd13603: log10_cal = 16'b0000010001111110;
            15'd13604: log10_cal = 16'b0000010001111110;
            15'd13605: log10_cal = 16'b0000010001111110;
            15'd13606: log10_cal = 16'b0000010001111110;
            15'd13607: log10_cal = 16'b0000010001111110;
            15'd13608: log10_cal = 16'b0000010001111110;
            15'd13609: log10_cal = 16'b0000010001111110;
            15'd13610: log10_cal = 16'b0000010001111110;
            15'd13611: log10_cal = 16'b0000010001111110;
            15'd13612: log10_cal = 16'b0000010001111110;
            15'd13613: log10_cal = 16'b0000010001111110;
            15'd13614: log10_cal = 16'b0000010001111110;
            15'd13615: log10_cal = 16'b0000010001111110;
            15'd13616: log10_cal = 16'b0000010001111110;
            15'd13617: log10_cal = 16'b0000010001111110;
            15'd13618: log10_cal = 16'b0000010001111110;
            15'd13619: log10_cal = 16'b0000010001111110;
            15'd13620: log10_cal = 16'b0000010001111110;
            15'd13621: log10_cal = 16'b0000010001111110;
            15'd13622: log10_cal = 16'b0000010001111110;
            15'd13623: log10_cal = 16'b0000010001111110;
            15'd13624: log10_cal = 16'b0000010001111110;
            15'd13625: log10_cal = 16'b0000010001111111;
            15'd13626: log10_cal = 16'b0000010001111111;
            15'd13627: log10_cal = 16'b0000010001111111;
            15'd13628: log10_cal = 16'b0000010001111111;
            15'd13629: log10_cal = 16'b0000010001111111;
            15'd13630: log10_cal = 16'b0000010001111111;
            15'd13631: log10_cal = 16'b0000010001111111;
            15'd13632: log10_cal = 16'b0000010001111111;
            15'd13633: log10_cal = 16'b0000010001111111;
            15'd13634: log10_cal = 16'b0000010001111111;
            15'd13635: log10_cal = 16'b0000010001111111;
            15'd13636: log10_cal = 16'b0000010001111111;
            15'd13637: log10_cal = 16'b0000010001111111;
            15'd13638: log10_cal = 16'b0000010001111111;
            15'd13639: log10_cal = 16'b0000010001111111;
            15'd13640: log10_cal = 16'b0000010001111111;
            15'd13641: log10_cal = 16'b0000010001111111;
            15'd13642: log10_cal = 16'b0000010001111111;
            15'd13643: log10_cal = 16'b0000010001111111;
            15'd13644: log10_cal = 16'b0000010001111111;
            15'd13645: log10_cal = 16'b0000010001111111;
            15'd13646: log10_cal = 16'b0000010001111111;
            15'd13647: log10_cal = 16'b0000010001111111;
            15'd13648: log10_cal = 16'b0000010001111111;
            15'd13649: log10_cal = 16'b0000010001111111;
            15'd13650: log10_cal = 16'b0000010001111111;
            15'd13651: log10_cal = 16'b0000010001111111;
            15'd13652: log10_cal = 16'b0000010001111111;
            15'd13653: log10_cal = 16'b0000010001111111;
            15'd13654: log10_cal = 16'b0000010001111111;
            15'd13655: log10_cal = 16'b0000010001111111;
            15'd13656: log10_cal = 16'b0000010010000000;
            15'd13657: log10_cal = 16'b0000010010000000;
            15'd13658: log10_cal = 16'b0000010010000000;
            15'd13659: log10_cal = 16'b0000010010000000;
            15'd13660: log10_cal = 16'b0000010010000000;
            15'd13661: log10_cal = 16'b0000010010000000;
            15'd13662: log10_cal = 16'b0000010010000000;
            15'd13663: log10_cal = 16'b0000010010000000;
            15'd13664: log10_cal = 16'b0000010010000000;
            15'd13665: log10_cal = 16'b0000010010000000;
            15'd13666: log10_cal = 16'b0000010010000000;
            15'd13667: log10_cal = 16'b0000010010000000;
            15'd13668: log10_cal = 16'b0000010010000000;
            15'd13669: log10_cal = 16'b0000010010000000;
            15'd13670: log10_cal = 16'b0000010010000000;
            15'd13671: log10_cal = 16'b0000010010000000;
            15'd13672: log10_cal = 16'b0000010010000000;
            15'd13673: log10_cal = 16'b0000010010000000;
            15'd13674: log10_cal = 16'b0000010010000000;
            15'd13675: log10_cal = 16'b0000010010000000;
            15'd13676: log10_cal = 16'b0000010010000000;
            15'd13677: log10_cal = 16'b0000010010000000;
            15'd13678: log10_cal = 16'b0000010010000000;
            15'd13679: log10_cal = 16'b0000010010000000;
            15'd13680: log10_cal = 16'b0000010010000000;
            15'd13681: log10_cal = 16'b0000010010000000;
            15'd13682: log10_cal = 16'b0000010010000000;
            15'd13683: log10_cal = 16'b0000010010000000;
            15'd13684: log10_cal = 16'b0000010010000000;
            15'd13685: log10_cal = 16'b0000010010000000;
            15'd13686: log10_cal = 16'b0000010010000001;
            15'd13687: log10_cal = 16'b0000010010000001;
            15'd13688: log10_cal = 16'b0000010010000001;
            15'd13689: log10_cal = 16'b0000010010000001;
            15'd13690: log10_cal = 16'b0000010010000001;
            15'd13691: log10_cal = 16'b0000010010000001;
            15'd13692: log10_cal = 16'b0000010010000001;
            15'd13693: log10_cal = 16'b0000010010000001;
            15'd13694: log10_cal = 16'b0000010010000001;
            15'd13695: log10_cal = 16'b0000010010000001;
            15'd13696: log10_cal = 16'b0000010010000001;
            15'd13697: log10_cal = 16'b0000010010000001;
            15'd13698: log10_cal = 16'b0000010010000001;
            15'd13699: log10_cal = 16'b0000010010000001;
            15'd13700: log10_cal = 16'b0000010010000001;
            15'd13701: log10_cal = 16'b0000010010000001;
            15'd13702: log10_cal = 16'b0000010010000001;
            15'd13703: log10_cal = 16'b0000010010000001;
            15'd13704: log10_cal = 16'b0000010010000001;
            15'd13705: log10_cal = 16'b0000010010000001;
            15'd13706: log10_cal = 16'b0000010010000001;
            15'd13707: log10_cal = 16'b0000010010000001;
            15'd13708: log10_cal = 16'b0000010010000001;
            15'd13709: log10_cal = 16'b0000010010000001;
            15'd13710: log10_cal = 16'b0000010010000001;
            15'd13711: log10_cal = 16'b0000010010000001;
            15'd13712: log10_cal = 16'b0000010010000001;
            15'd13713: log10_cal = 16'b0000010010000001;
            15'd13714: log10_cal = 16'b0000010010000001;
            15'd13715: log10_cal = 16'b0000010010000001;
            15'd13716: log10_cal = 16'b0000010010000001;
            15'd13717: log10_cal = 16'b0000010010000010;
            15'd13718: log10_cal = 16'b0000010010000010;
            15'd13719: log10_cal = 16'b0000010010000010;
            15'd13720: log10_cal = 16'b0000010010000010;
            15'd13721: log10_cal = 16'b0000010010000010;
            15'd13722: log10_cal = 16'b0000010010000010;
            15'd13723: log10_cal = 16'b0000010010000010;
            15'd13724: log10_cal = 16'b0000010010000010;
            15'd13725: log10_cal = 16'b0000010010000010;
            15'd13726: log10_cal = 16'b0000010010000010;
            15'd13727: log10_cal = 16'b0000010010000010;
            15'd13728: log10_cal = 16'b0000010010000010;
            15'd13729: log10_cal = 16'b0000010010000010;
            15'd13730: log10_cal = 16'b0000010010000010;
            15'd13731: log10_cal = 16'b0000010010000010;
            15'd13732: log10_cal = 16'b0000010010000010;
            15'd13733: log10_cal = 16'b0000010010000010;
            15'd13734: log10_cal = 16'b0000010010000010;
            15'd13735: log10_cal = 16'b0000010010000010;
            15'd13736: log10_cal = 16'b0000010010000010;
            15'd13737: log10_cal = 16'b0000010010000010;
            15'd13738: log10_cal = 16'b0000010010000010;
            15'd13739: log10_cal = 16'b0000010010000010;
            15'd13740: log10_cal = 16'b0000010010000010;
            15'd13741: log10_cal = 16'b0000010010000010;
            15'd13742: log10_cal = 16'b0000010010000010;
            15'd13743: log10_cal = 16'b0000010010000010;
            15'd13744: log10_cal = 16'b0000010010000010;
            15'd13745: log10_cal = 16'b0000010010000010;
            15'd13746: log10_cal = 16'b0000010010000010;
            15'd13747: log10_cal = 16'b0000010010000010;
            15'd13748: log10_cal = 16'b0000010010000011;
            15'd13749: log10_cal = 16'b0000010010000011;
            15'd13750: log10_cal = 16'b0000010010000011;
            15'd13751: log10_cal = 16'b0000010010000011;
            15'd13752: log10_cal = 16'b0000010010000011;
            15'd13753: log10_cal = 16'b0000010010000011;
            15'd13754: log10_cal = 16'b0000010010000011;
            15'd13755: log10_cal = 16'b0000010010000011;
            15'd13756: log10_cal = 16'b0000010010000011;
            15'd13757: log10_cal = 16'b0000010010000011;
            15'd13758: log10_cal = 16'b0000010010000011;
            15'd13759: log10_cal = 16'b0000010010000011;
            15'd13760: log10_cal = 16'b0000010010000011;
            15'd13761: log10_cal = 16'b0000010010000011;
            15'd13762: log10_cal = 16'b0000010010000011;
            15'd13763: log10_cal = 16'b0000010010000011;
            15'd13764: log10_cal = 16'b0000010010000011;
            15'd13765: log10_cal = 16'b0000010010000011;
            15'd13766: log10_cal = 16'b0000010010000011;
            15'd13767: log10_cal = 16'b0000010010000011;
            15'd13768: log10_cal = 16'b0000010010000011;
            15'd13769: log10_cal = 16'b0000010010000011;
            15'd13770: log10_cal = 16'b0000010010000011;
            15'd13771: log10_cal = 16'b0000010010000011;
            15'd13772: log10_cal = 16'b0000010010000011;
            15'd13773: log10_cal = 16'b0000010010000011;
            15'd13774: log10_cal = 16'b0000010010000011;
            15'd13775: log10_cal = 16'b0000010010000011;
            15'd13776: log10_cal = 16'b0000010010000011;
            15'd13777: log10_cal = 16'b0000010010000011;
            15'd13778: log10_cal = 16'b0000010010000011;
            15'd13779: log10_cal = 16'b0000010010000100;
            15'd13780: log10_cal = 16'b0000010010000100;
            15'd13781: log10_cal = 16'b0000010010000100;
            15'd13782: log10_cal = 16'b0000010010000100;
            15'd13783: log10_cal = 16'b0000010010000100;
            15'd13784: log10_cal = 16'b0000010010000100;
            15'd13785: log10_cal = 16'b0000010010000100;
            15'd13786: log10_cal = 16'b0000010010000100;
            15'd13787: log10_cal = 16'b0000010010000100;
            15'd13788: log10_cal = 16'b0000010010000100;
            15'd13789: log10_cal = 16'b0000010010000100;
            15'd13790: log10_cal = 16'b0000010010000100;
            15'd13791: log10_cal = 16'b0000010010000100;
            15'd13792: log10_cal = 16'b0000010010000100;
            15'd13793: log10_cal = 16'b0000010010000100;
            15'd13794: log10_cal = 16'b0000010010000100;
            15'd13795: log10_cal = 16'b0000010010000100;
            15'd13796: log10_cal = 16'b0000010010000100;
            15'd13797: log10_cal = 16'b0000010010000100;
            15'd13798: log10_cal = 16'b0000010010000100;
            15'd13799: log10_cal = 16'b0000010010000100;
            15'd13800: log10_cal = 16'b0000010010000100;
            15'd13801: log10_cal = 16'b0000010010000100;
            15'd13802: log10_cal = 16'b0000010010000100;
            15'd13803: log10_cal = 16'b0000010010000100;
            15'd13804: log10_cal = 16'b0000010010000100;
            15'd13805: log10_cal = 16'b0000010010000100;
            15'd13806: log10_cal = 16'b0000010010000100;
            15'd13807: log10_cal = 16'b0000010010000100;
            15'd13808: log10_cal = 16'b0000010010000100;
            15'd13809: log10_cal = 16'b0000010010000100;
            15'd13810: log10_cal = 16'b0000010010000101;
            15'd13811: log10_cal = 16'b0000010010000101;
            15'd13812: log10_cal = 16'b0000010010000101;
            15'd13813: log10_cal = 16'b0000010010000101;
            15'd13814: log10_cal = 16'b0000010010000101;
            15'd13815: log10_cal = 16'b0000010010000101;
            15'd13816: log10_cal = 16'b0000010010000101;
            15'd13817: log10_cal = 16'b0000010010000101;
            15'd13818: log10_cal = 16'b0000010010000101;
            15'd13819: log10_cal = 16'b0000010010000101;
            15'd13820: log10_cal = 16'b0000010010000101;
            15'd13821: log10_cal = 16'b0000010010000101;
            15'd13822: log10_cal = 16'b0000010010000101;
            15'd13823: log10_cal = 16'b0000010010000101;
            15'd13824: log10_cal = 16'b0000010010000101;
            15'd13825: log10_cal = 16'b0000010010000101;
            15'd13826: log10_cal = 16'b0000010010000101;
            15'd13827: log10_cal = 16'b0000010010000101;
            15'd13828: log10_cal = 16'b0000010010000101;
            15'd13829: log10_cal = 16'b0000010010000101;
            15'd13830: log10_cal = 16'b0000010010000101;
            15'd13831: log10_cal = 16'b0000010010000101;
            15'd13832: log10_cal = 16'b0000010010000101;
            15'd13833: log10_cal = 16'b0000010010000101;
            15'd13834: log10_cal = 16'b0000010010000101;
            15'd13835: log10_cal = 16'b0000010010000101;
            15'd13836: log10_cal = 16'b0000010010000101;
            15'd13837: log10_cal = 16'b0000010010000101;
            15'd13838: log10_cal = 16'b0000010010000101;
            15'd13839: log10_cal = 16'b0000010010000101;
            15'd13840: log10_cal = 16'b0000010010000101;
            15'd13841: log10_cal = 16'b0000010010000110;
            15'd13842: log10_cal = 16'b0000010010000110;
            15'd13843: log10_cal = 16'b0000010010000110;
            15'd13844: log10_cal = 16'b0000010010000110;
            15'd13845: log10_cal = 16'b0000010010000110;
            15'd13846: log10_cal = 16'b0000010010000110;
            15'd13847: log10_cal = 16'b0000010010000110;
            15'd13848: log10_cal = 16'b0000010010000110;
            15'd13849: log10_cal = 16'b0000010010000110;
            15'd13850: log10_cal = 16'b0000010010000110;
            15'd13851: log10_cal = 16'b0000010010000110;
            15'd13852: log10_cal = 16'b0000010010000110;
            15'd13853: log10_cal = 16'b0000010010000110;
            15'd13854: log10_cal = 16'b0000010010000110;
            15'd13855: log10_cal = 16'b0000010010000110;
            15'd13856: log10_cal = 16'b0000010010000110;
            15'd13857: log10_cal = 16'b0000010010000110;
            15'd13858: log10_cal = 16'b0000010010000110;
            15'd13859: log10_cal = 16'b0000010010000110;
            15'd13860: log10_cal = 16'b0000010010000110;
            15'd13861: log10_cal = 16'b0000010010000110;
            15'd13862: log10_cal = 16'b0000010010000110;
            15'd13863: log10_cal = 16'b0000010010000110;
            15'd13864: log10_cal = 16'b0000010010000110;
            15'd13865: log10_cal = 16'b0000010010000110;
            15'd13866: log10_cal = 16'b0000010010000110;
            15'd13867: log10_cal = 16'b0000010010000110;
            15'd13868: log10_cal = 16'b0000010010000110;
            15'd13869: log10_cal = 16'b0000010010000110;
            15'd13870: log10_cal = 16'b0000010010000110;
            15'd13871: log10_cal = 16'b0000010010000110;
            15'd13872: log10_cal = 16'b0000010010000111;
            15'd13873: log10_cal = 16'b0000010010000111;
            15'd13874: log10_cal = 16'b0000010010000111;
            15'd13875: log10_cal = 16'b0000010010000111;
            15'd13876: log10_cal = 16'b0000010010000111;
            15'd13877: log10_cal = 16'b0000010010000111;
            15'd13878: log10_cal = 16'b0000010010000111;
            15'd13879: log10_cal = 16'b0000010010000111;
            15'd13880: log10_cal = 16'b0000010010000111;
            15'd13881: log10_cal = 16'b0000010010000111;
            15'd13882: log10_cal = 16'b0000010010000111;
            15'd13883: log10_cal = 16'b0000010010000111;
            15'd13884: log10_cal = 16'b0000010010000111;
            15'd13885: log10_cal = 16'b0000010010000111;
            15'd13886: log10_cal = 16'b0000010010000111;
            15'd13887: log10_cal = 16'b0000010010000111;
            15'd13888: log10_cal = 16'b0000010010000111;
            15'd13889: log10_cal = 16'b0000010010000111;
            15'd13890: log10_cal = 16'b0000010010000111;
            15'd13891: log10_cal = 16'b0000010010000111;
            15'd13892: log10_cal = 16'b0000010010000111;
            15'd13893: log10_cal = 16'b0000010010000111;
            15'd13894: log10_cal = 16'b0000010010000111;
            15'd13895: log10_cal = 16'b0000010010000111;
            15'd13896: log10_cal = 16'b0000010010000111;
            15'd13897: log10_cal = 16'b0000010010000111;
            15'd13898: log10_cal = 16'b0000010010000111;
            15'd13899: log10_cal = 16'b0000010010000111;
            15'd13900: log10_cal = 16'b0000010010000111;
            15'd13901: log10_cal = 16'b0000010010000111;
            15'd13902: log10_cal = 16'b0000010010000111;
            15'd13903: log10_cal = 16'b0000010010000111;
            15'd13904: log10_cal = 16'b0000010010001000;
            15'd13905: log10_cal = 16'b0000010010001000;
            15'd13906: log10_cal = 16'b0000010010001000;
            15'd13907: log10_cal = 16'b0000010010001000;
            15'd13908: log10_cal = 16'b0000010010001000;
            15'd13909: log10_cal = 16'b0000010010001000;
            15'd13910: log10_cal = 16'b0000010010001000;
            15'd13911: log10_cal = 16'b0000010010001000;
            15'd13912: log10_cal = 16'b0000010010001000;
            15'd13913: log10_cal = 16'b0000010010001000;
            15'd13914: log10_cal = 16'b0000010010001000;
            15'd13915: log10_cal = 16'b0000010010001000;
            15'd13916: log10_cal = 16'b0000010010001000;
            15'd13917: log10_cal = 16'b0000010010001000;
            15'd13918: log10_cal = 16'b0000010010001000;
            15'd13919: log10_cal = 16'b0000010010001000;
            15'd13920: log10_cal = 16'b0000010010001000;
            15'd13921: log10_cal = 16'b0000010010001000;
            15'd13922: log10_cal = 16'b0000010010001000;
            15'd13923: log10_cal = 16'b0000010010001000;
            15'd13924: log10_cal = 16'b0000010010001000;
            15'd13925: log10_cal = 16'b0000010010001000;
            15'd13926: log10_cal = 16'b0000010010001000;
            15'd13927: log10_cal = 16'b0000010010001000;
            15'd13928: log10_cal = 16'b0000010010001000;
            15'd13929: log10_cal = 16'b0000010010001000;
            15'd13930: log10_cal = 16'b0000010010001000;
            15'd13931: log10_cal = 16'b0000010010001000;
            15'd13932: log10_cal = 16'b0000010010001000;
            15'd13933: log10_cal = 16'b0000010010001000;
            15'd13934: log10_cal = 16'b0000010010001000;
            15'd13935: log10_cal = 16'b0000010010001001;
            15'd13936: log10_cal = 16'b0000010010001001;
            15'd13937: log10_cal = 16'b0000010010001001;
            15'd13938: log10_cal = 16'b0000010010001001;
            15'd13939: log10_cal = 16'b0000010010001001;
            15'd13940: log10_cal = 16'b0000010010001001;
            15'd13941: log10_cal = 16'b0000010010001001;
            15'd13942: log10_cal = 16'b0000010010001001;
            15'd13943: log10_cal = 16'b0000010010001001;
            15'd13944: log10_cal = 16'b0000010010001001;
            15'd13945: log10_cal = 16'b0000010010001001;
            15'd13946: log10_cal = 16'b0000010010001001;
            15'd13947: log10_cal = 16'b0000010010001001;
            15'd13948: log10_cal = 16'b0000010010001001;
            15'd13949: log10_cal = 16'b0000010010001001;
            15'd13950: log10_cal = 16'b0000010010001001;
            15'd13951: log10_cal = 16'b0000010010001001;
            15'd13952: log10_cal = 16'b0000010010001001;
            15'd13953: log10_cal = 16'b0000010010001001;
            15'd13954: log10_cal = 16'b0000010010001001;
            15'd13955: log10_cal = 16'b0000010010001001;
            15'd13956: log10_cal = 16'b0000010010001001;
            15'd13957: log10_cal = 16'b0000010010001001;
            15'd13958: log10_cal = 16'b0000010010001001;
            15'd13959: log10_cal = 16'b0000010010001001;
            15'd13960: log10_cal = 16'b0000010010001001;
            15'd13961: log10_cal = 16'b0000010010001001;
            15'd13962: log10_cal = 16'b0000010010001001;
            15'd13963: log10_cal = 16'b0000010010001001;
            15'd13964: log10_cal = 16'b0000010010001001;
            15'd13965: log10_cal = 16'b0000010010001001;
            15'd13966: log10_cal = 16'b0000010010001010;
            15'd13967: log10_cal = 16'b0000010010001010;
            15'd13968: log10_cal = 16'b0000010010001010;
            15'd13969: log10_cal = 16'b0000010010001010;
            15'd13970: log10_cal = 16'b0000010010001010;
            15'd13971: log10_cal = 16'b0000010010001010;
            15'd13972: log10_cal = 16'b0000010010001010;
            15'd13973: log10_cal = 16'b0000010010001010;
            15'd13974: log10_cal = 16'b0000010010001010;
            15'd13975: log10_cal = 16'b0000010010001010;
            15'd13976: log10_cal = 16'b0000010010001010;
            15'd13977: log10_cal = 16'b0000010010001010;
            15'd13978: log10_cal = 16'b0000010010001010;
            15'd13979: log10_cal = 16'b0000010010001010;
            15'd13980: log10_cal = 16'b0000010010001010;
            15'd13981: log10_cal = 16'b0000010010001010;
            15'd13982: log10_cal = 16'b0000010010001010;
            15'd13983: log10_cal = 16'b0000010010001010;
            15'd13984: log10_cal = 16'b0000010010001010;
            15'd13985: log10_cal = 16'b0000010010001010;
            15'd13986: log10_cal = 16'b0000010010001010;
            15'd13987: log10_cal = 16'b0000010010001010;
            15'd13988: log10_cal = 16'b0000010010001010;
            15'd13989: log10_cal = 16'b0000010010001010;
            15'd13990: log10_cal = 16'b0000010010001010;
            15'd13991: log10_cal = 16'b0000010010001010;
            15'd13992: log10_cal = 16'b0000010010001010;
            15'd13993: log10_cal = 16'b0000010010001010;
            15'd13994: log10_cal = 16'b0000010010001010;
            15'd13995: log10_cal = 16'b0000010010001010;
            15'd13996: log10_cal = 16'b0000010010001010;
            15'd13997: log10_cal = 16'b0000010010001010;
            15'd13998: log10_cal = 16'b0000010010001011;
            15'd13999: log10_cal = 16'b0000010010001011;
            15'd14000: log10_cal = 16'b0000010010001011;
            15'd14001: log10_cal = 16'b0000010010001011;
            15'd14002: log10_cal = 16'b0000010010001011;
            15'd14003: log10_cal = 16'b0000010010001011;
            15'd14004: log10_cal = 16'b0000010010001011;
            15'd14005: log10_cal = 16'b0000010010001011;
            15'd14006: log10_cal = 16'b0000010010001011;
            15'd14007: log10_cal = 16'b0000010010001011;
            15'd14008: log10_cal = 16'b0000010010001011;
            15'd14009: log10_cal = 16'b0000010010001011;
            15'd14010: log10_cal = 16'b0000010010001011;
            15'd14011: log10_cal = 16'b0000010010001011;
            15'd14012: log10_cal = 16'b0000010010001011;
            15'd14013: log10_cal = 16'b0000010010001011;
            15'd14014: log10_cal = 16'b0000010010001011;
            15'd14015: log10_cal = 16'b0000010010001011;
            15'd14016: log10_cal = 16'b0000010010001011;
            15'd14017: log10_cal = 16'b0000010010001011;
            15'd14018: log10_cal = 16'b0000010010001011;
            15'd14019: log10_cal = 16'b0000010010001011;
            15'd14020: log10_cal = 16'b0000010010001011;
            15'd14021: log10_cal = 16'b0000010010001011;
            15'd14022: log10_cal = 16'b0000010010001011;
            15'd14023: log10_cal = 16'b0000010010001011;
            15'd14024: log10_cal = 16'b0000010010001011;
            15'd14025: log10_cal = 16'b0000010010001011;
            15'd14026: log10_cal = 16'b0000010010001011;
            15'd14027: log10_cal = 16'b0000010010001011;
            15'd14028: log10_cal = 16'b0000010010001011;
            15'd14029: log10_cal = 16'b0000010010001100;
            15'd14030: log10_cal = 16'b0000010010001100;
            15'd14031: log10_cal = 16'b0000010010001100;
            15'd14032: log10_cal = 16'b0000010010001100;
            15'd14033: log10_cal = 16'b0000010010001100;
            15'd14034: log10_cal = 16'b0000010010001100;
            15'd14035: log10_cal = 16'b0000010010001100;
            15'd14036: log10_cal = 16'b0000010010001100;
            15'd14037: log10_cal = 16'b0000010010001100;
            15'd14038: log10_cal = 16'b0000010010001100;
            15'd14039: log10_cal = 16'b0000010010001100;
            15'd14040: log10_cal = 16'b0000010010001100;
            15'd14041: log10_cal = 16'b0000010010001100;
            15'd14042: log10_cal = 16'b0000010010001100;
            15'd14043: log10_cal = 16'b0000010010001100;
            15'd14044: log10_cal = 16'b0000010010001100;
            15'd14045: log10_cal = 16'b0000010010001100;
            15'd14046: log10_cal = 16'b0000010010001100;
            15'd14047: log10_cal = 16'b0000010010001100;
            15'd14048: log10_cal = 16'b0000010010001100;
            15'd14049: log10_cal = 16'b0000010010001100;
            15'd14050: log10_cal = 16'b0000010010001100;
            15'd14051: log10_cal = 16'b0000010010001100;
            15'd14052: log10_cal = 16'b0000010010001100;
            15'd14053: log10_cal = 16'b0000010010001100;
            15'd14054: log10_cal = 16'b0000010010001100;
            15'd14055: log10_cal = 16'b0000010010001100;
            15'd14056: log10_cal = 16'b0000010010001100;
            15'd14057: log10_cal = 16'b0000010010001100;
            15'd14058: log10_cal = 16'b0000010010001100;
            15'd14059: log10_cal = 16'b0000010010001100;
            15'd14060: log10_cal = 16'b0000010010001100;
            15'd14061: log10_cal = 16'b0000010010001101;
            15'd14062: log10_cal = 16'b0000010010001101;
            15'd14063: log10_cal = 16'b0000010010001101;
            15'd14064: log10_cal = 16'b0000010010001101;
            15'd14065: log10_cal = 16'b0000010010001101;
            15'd14066: log10_cal = 16'b0000010010001101;
            15'd14067: log10_cal = 16'b0000010010001101;
            15'd14068: log10_cal = 16'b0000010010001101;
            15'd14069: log10_cal = 16'b0000010010001101;
            15'd14070: log10_cal = 16'b0000010010001101;
            15'd14071: log10_cal = 16'b0000010010001101;
            15'd14072: log10_cal = 16'b0000010010001101;
            15'd14073: log10_cal = 16'b0000010010001101;
            15'd14074: log10_cal = 16'b0000010010001101;
            15'd14075: log10_cal = 16'b0000010010001101;
            15'd14076: log10_cal = 16'b0000010010001101;
            15'd14077: log10_cal = 16'b0000010010001101;
            15'd14078: log10_cal = 16'b0000010010001101;
            15'd14079: log10_cal = 16'b0000010010001101;
            15'd14080: log10_cal = 16'b0000010010001101;
            15'd14081: log10_cal = 16'b0000010010001101;
            15'd14082: log10_cal = 16'b0000010010001101;
            15'd14083: log10_cal = 16'b0000010010001101;
            15'd14084: log10_cal = 16'b0000010010001101;
            15'd14085: log10_cal = 16'b0000010010001101;
            15'd14086: log10_cal = 16'b0000010010001101;
            15'd14087: log10_cal = 16'b0000010010001101;
            15'd14088: log10_cal = 16'b0000010010001101;
            15'd14089: log10_cal = 16'b0000010010001101;
            15'd14090: log10_cal = 16'b0000010010001101;
            15'd14091: log10_cal = 16'b0000010010001101;
            15'd14092: log10_cal = 16'b0000010010001110;
            15'd14093: log10_cal = 16'b0000010010001110;
            15'd14094: log10_cal = 16'b0000010010001110;
            15'd14095: log10_cal = 16'b0000010010001110;
            15'd14096: log10_cal = 16'b0000010010001110;
            15'd14097: log10_cal = 16'b0000010010001110;
            15'd14098: log10_cal = 16'b0000010010001110;
            15'd14099: log10_cal = 16'b0000010010001110;
            15'd14100: log10_cal = 16'b0000010010001110;
            15'd14101: log10_cal = 16'b0000010010001110;
            15'd14102: log10_cal = 16'b0000010010001110;
            15'd14103: log10_cal = 16'b0000010010001110;
            15'd14104: log10_cal = 16'b0000010010001110;
            15'd14105: log10_cal = 16'b0000010010001110;
            15'd14106: log10_cal = 16'b0000010010001110;
            15'd14107: log10_cal = 16'b0000010010001110;
            15'd14108: log10_cal = 16'b0000010010001110;
            15'd14109: log10_cal = 16'b0000010010001110;
            15'd14110: log10_cal = 16'b0000010010001110;
            15'd14111: log10_cal = 16'b0000010010001110;
            15'd14112: log10_cal = 16'b0000010010001110;
            15'd14113: log10_cal = 16'b0000010010001110;
            15'd14114: log10_cal = 16'b0000010010001110;
            15'd14115: log10_cal = 16'b0000010010001110;
            15'd14116: log10_cal = 16'b0000010010001110;
            15'd14117: log10_cal = 16'b0000010010001110;
            15'd14118: log10_cal = 16'b0000010010001110;
            15'd14119: log10_cal = 16'b0000010010001110;
            15'd14120: log10_cal = 16'b0000010010001110;
            15'd14121: log10_cal = 16'b0000010010001110;
            15'd14122: log10_cal = 16'b0000010010001110;
            15'd14123: log10_cal = 16'b0000010010001110;
            15'd14124: log10_cal = 16'b0000010010001111;
            15'd14125: log10_cal = 16'b0000010010001111;
            15'd14126: log10_cal = 16'b0000010010001111;
            15'd14127: log10_cal = 16'b0000010010001111;
            15'd14128: log10_cal = 16'b0000010010001111;
            15'd14129: log10_cal = 16'b0000010010001111;
            15'd14130: log10_cal = 16'b0000010010001111;
            15'd14131: log10_cal = 16'b0000010010001111;
            15'd14132: log10_cal = 16'b0000010010001111;
            15'd14133: log10_cal = 16'b0000010010001111;
            15'd14134: log10_cal = 16'b0000010010001111;
            15'd14135: log10_cal = 16'b0000010010001111;
            15'd14136: log10_cal = 16'b0000010010001111;
            15'd14137: log10_cal = 16'b0000010010001111;
            15'd14138: log10_cal = 16'b0000010010001111;
            15'd14139: log10_cal = 16'b0000010010001111;
            15'd14140: log10_cal = 16'b0000010010001111;
            15'd14141: log10_cal = 16'b0000010010001111;
            15'd14142: log10_cal = 16'b0000010010001111;
            15'd14143: log10_cal = 16'b0000010010001111;
            15'd14144: log10_cal = 16'b0000010010001111;
            15'd14145: log10_cal = 16'b0000010010001111;
            15'd14146: log10_cal = 16'b0000010010001111;
            15'd14147: log10_cal = 16'b0000010010001111;
            15'd14148: log10_cal = 16'b0000010010001111;
            15'd14149: log10_cal = 16'b0000010010001111;
            15'd14150: log10_cal = 16'b0000010010001111;
            15'd14151: log10_cal = 16'b0000010010001111;
            15'd14152: log10_cal = 16'b0000010010001111;
            15'd14153: log10_cal = 16'b0000010010001111;
            15'd14154: log10_cal = 16'b0000010010001111;
            15'd14155: log10_cal = 16'b0000010010001111;
            15'd14156: log10_cal = 16'b0000010010010000;
            15'd14157: log10_cal = 16'b0000010010010000;
            15'd14158: log10_cal = 16'b0000010010010000;
            15'd14159: log10_cal = 16'b0000010010010000;
            15'd14160: log10_cal = 16'b0000010010010000;
            15'd14161: log10_cal = 16'b0000010010010000;
            15'd14162: log10_cal = 16'b0000010010010000;
            15'd14163: log10_cal = 16'b0000010010010000;
            15'd14164: log10_cal = 16'b0000010010010000;
            15'd14165: log10_cal = 16'b0000010010010000;
            15'd14166: log10_cal = 16'b0000010010010000;
            15'd14167: log10_cal = 16'b0000010010010000;
            15'd14168: log10_cal = 16'b0000010010010000;
            15'd14169: log10_cal = 16'b0000010010010000;
            15'd14170: log10_cal = 16'b0000010010010000;
            15'd14171: log10_cal = 16'b0000010010010000;
            15'd14172: log10_cal = 16'b0000010010010000;
            15'd14173: log10_cal = 16'b0000010010010000;
            15'd14174: log10_cal = 16'b0000010010010000;
            15'd14175: log10_cal = 16'b0000010010010000;
            15'd14176: log10_cal = 16'b0000010010010000;
            15'd14177: log10_cal = 16'b0000010010010000;
            15'd14178: log10_cal = 16'b0000010010010000;
            15'd14179: log10_cal = 16'b0000010010010000;
            15'd14180: log10_cal = 16'b0000010010010000;
            15'd14181: log10_cal = 16'b0000010010010000;
            15'd14182: log10_cal = 16'b0000010010010000;
            15'd14183: log10_cal = 16'b0000010010010000;
            15'd14184: log10_cal = 16'b0000010010010000;
            15'd14185: log10_cal = 16'b0000010010010000;
            15'd14186: log10_cal = 16'b0000010010010000;
            15'd14187: log10_cal = 16'b0000010010010000;
            15'd14188: log10_cal = 16'b0000010010010001;
            15'd14189: log10_cal = 16'b0000010010010001;
            15'd14190: log10_cal = 16'b0000010010010001;
            15'd14191: log10_cal = 16'b0000010010010001;
            15'd14192: log10_cal = 16'b0000010010010001;
            15'd14193: log10_cal = 16'b0000010010010001;
            15'd14194: log10_cal = 16'b0000010010010001;
            15'd14195: log10_cal = 16'b0000010010010001;
            15'd14196: log10_cal = 16'b0000010010010001;
            15'd14197: log10_cal = 16'b0000010010010001;
            15'd14198: log10_cal = 16'b0000010010010001;
            15'd14199: log10_cal = 16'b0000010010010001;
            15'd14200: log10_cal = 16'b0000010010010001;
            15'd14201: log10_cal = 16'b0000010010010001;
            15'd14202: log10_cal = 16'b0000010010010001;
            15'd14203: log10_cal = 16'b0000010010010001;
            15'd14204: log10_cal = 16'b0000010010010001;
            15'd14205: log10_cal = 16'b0000010010010001;
            15'd14206: log10_cal = 16'b0000010010010001;
            15'd14207: log10_cal = 16'b0000010010010001;
            15'd14208: log10_cal = 16'b0000010010010001;
            15'd14209: log10_cal = 16'b0000010010010001;
            15'd14210: log10_cal = 16'b0000010010010001;
            15'd14211: log10_cal = 16'b0000010010010001;
            15'd14212: log10_cal = 16'b0000010010010001;
            15'd14213: log10_cal = 16'b0000010010010001;
            15'd14214: log10_cal = 16'b0000010010010001;
            15'd14215: log10_cal = 16'b0000010010010001;
            15'd14216: log10_cal = 16'b0000010010010001;
            15'd14217: log10_cal = 16'b0000010010010001;
            15'd14218: log10_cal = 16'b0000010010010001;
            15'd14219: log10_cal = 16'b0000010010010001;
            15'd14220: log10_cal = 16'b0000010010010010;
            15'd14221: log10_cal = 16'b0000010010010010;
            15'd14222: log10_cal = 16'b0000010010010010;
            15'd14223: log10_cal = 16'b0000010010010010;
            15'd14224: log10_cal = 16'b0000010010010010;
            15'd14225: log10_cal = 16'b0000010010010010;
            15'd14226: log10_cal = 16'b0000010010010010;
            15'd14227: log10_cal = 16'b0000010010010010;
            15'd14228: log10_cal = 16'b0000010010010010;
            15'd14229: log10_cal = 16'b0000010010010010;
            15'd14230: log10_cal = 16'b0000010010010010;
            15'd14231: log10_cal = 16'b0000010010010010;
            15'd14232: log10_cal = 16'b0000010010010010;
            15'd14233: log10_cal = 16'b0000010010010010;
            15'd14234: log10_cal = 16'b0000010010010010;
            15'd14235: log10_cal = 16'b0000010010010010;
            15'd14236: log10_cal = 16'b0000010010010010;
            15'd14237: log10_cal = 16'b0000010010010010;
            15'd14238: log10_cal = 16'b0000010010010010;
            15'd14239: log10_cal = 16'b0000010010010010;
            15'd14240: log10_cal = 16'b0000010010010010;
            15'd14241: log10_cal = 16'b0000010010010010;
            15'd14242: log10_cal = 16'b0000010010010010;
            15'd14243: log10_cal = 16'b0000010010010010;
            15'd14244: log10_cal = 16'b0000010010010010;
            15'd14245: log10_cal = 16'b0000010010010010;
            15'd14246: log10_cal = 16'b0000010010010010;
            15'd14247: log10_cal = 16'b0000010010010010;
            15'd14248: log10_cal = 16'b0000010010010010;
            15'd14249: log10_cal = 16'b0000010010010010;
            15'd14250: log10_cal = 16'b0000010010010010;
            15'd14251: log10_cal = 16'b0000010010010010;
            15'd14252: log10_cal = 16'b0000010010010011;
            15'd14253: log10_cal = 16'b0000010010010011;
            15'd14254: log10_cal = 16'b0000010010010011;
            15'd14255: log10_cal = 16'b0000010010010011;
            15'd14256: log10_cal = 16'b0000010010010011;
            15'd14257: log10_cal = 16'b0000010010010011;
            15'd14258: log10_cal = 16'b0000010010010011;
            15'd14259: log10_cal = 16'b0000010010010011;
            15'd14260: log10_cal = 16'b0000010010010011;
            15'd14261: log10_cal = 16'b0000010010010011;
            15'd14262: log10_cal = 16'b0000010010010011;
            15'd14263: log10_cal = 16'b0000010010010011;
            15'd14264: log10_cal = 16'b0000010010010011;
            15'd14265: log10_cal = 16'b0000010010010011;
            15'd14266: log10_cal = 16'b0000010010010011;
            15'd14267: log10_cal = 16'b0000010010010011;
            15'd14268: log10_cal = 16'b0000010010010011;
            15'd14269: log10_cal = 16'b0000010010010011;
            15'd14270: log10_cal = 16'b0000010010010011;
            15'd14271: log10_cal = 16'b0000010010010011;
            15'd14272: log10_cal = 16'b0000010010010011;
            15'd14273: log10_cal = 16'b0000010010010011;
            15'd14274: log10_cal = 16'b0000010010010011;
            15'd14275: log10_cal = 16'b0000010010010011;
            15'd14276: log10_cal = 16'b0000010010010011;
            15'd14277: log10_cal = 16'b0000010010010011;
            15'd14278: log10_cal = 16'b0000010010010011;
            15'd14279: log10_cal = 16'b0000010010010011;
            15'd14280: log10_cal = 16'b0000010010010011;
            15'd14281: log10_cal = 16'b0000010010010011;
            15'd14282: log10_cal = 16'b0000010010010011;
            15'd14283: log10_cal = 16'b0000010010010011;
            15'd14284: log10_cal = 16'b0000010010010100;
            15'd14285: log10_cal = 16'b0000010010010100;
            15'd14286: log10_cal = 16'b0000010010010100;
            15'd14287: log10_cal = 16'b0000010010010100;
            15'd14288: log10_cal = 16'b0000010010010100;
            15'd14289: log10_cal = 16'b0000010010010100;
            15'd14290: log10_cal = 16'b0000010010010100;
            15'd14291: log10_cal = 16'b0000010010010100;
            15'd14292: log10_cal = 16'b0000010010010100;
            15'd14293: log10_cal = 16'b0000010010010100;
            15'd14294: log10_cal = 16'b0000010010010100;
            15'd14295: log10_cal = 16'b0000010010010100;
            15'd14296: log10_cal = 16'b0000010010010100;
            15'd14297: log10_cal = 16'b0000010010010100;
            15'd14298: log10_cal = 16'b0000010010010100;
            15'd14299: log10_cal = 16'b0000010010010100;
            15'd14300: log10_cal = 16'b0000010010010100;
            15'd14301: log10_cal = 16'b0000010010010100;
            15'd14302: log10_cal = 16'b0000010010010100;
            15'd14303: log10_cal = 16'b0000010010010100;
            15'd14304: log10_cal = 16'b0000010010010100;
            15'd14305: log10_cal = 16'b0000010010010100;
            15'd14306: log10_cal = 16'b0000010010010100;
            15'd14307: log10_cal = 16'b0000010010010100;
            15'd14308: log10_cal = 16'b0000010010010100;
            15'd14309: log10_cal = 16'b0000010010010100;
            15'd14310: log10_cal = 16'b0000010010010100;
            15'd14311: log10_cal = 16'b0000010010010100;
            15'd14312: log10_cal = 16'b0000010010010100;
            15'd14313: log10_cal = 16'b0000010010010100;
            15'd14314: log10_cal = 16'b0000010010010100;
            15'd14315: log10_cal = 16'b0000010010010100;
            15'd14316: log10_cal = 16'b0000010010010101;
            15'd14317: log10_cal = 16'b0000010010010101;
            15'd14318: log10_cal = 16'b0000010010010101;
            15'd14319: log10_cal = 16'b0000010010010101;
            15'd14320: log10_cal = 16'b0000010010010101;
            15'd14321: log10_cal = 16'b0000010010010101;
            15'd14322: log10_cal = 16'b0000010010010101;
            15'd14323: log10_cal = 16'b0000010010010101;
            15'd14324: log10_cal = 16'b0000010010010101;
            15'd14325: log10_cal = 16'b0000010010010101;
            15'd14326: log10_cal = 16'b0000010010010101;
            15'd14327: log10_cal = 16'b0000010010010101;
            15'd14328: log10_cal = 16'b0000010010010101;
            15'd14329: log10_cal = 16'b0000010010010101;
            15'd14330: log10_cal = 16'b0000010010010101;
            15'd14331: log10_cal = 16'b0000010010010101;
            15'd14332: log10_cal = 16'b0000010010010101;
            15'd14333: log10_cal = 16'b0000010010010101;
            15'd14334: log10_cal = 16'b0000010010010101;
            15'd14335: log10_cal = 16'b0000010010010101;
            15'd14336: log10_cal = 16'b0000010010010101;
            15'd14337: log10_cal = 16'b0000010010010101;
            15'd14338: log10_cal = 16'b0000010010010101;
            15'd14339: log10_cal = 16'b0000010010010101;
            15'd14340: log10_cal = 16'b0000010010010101;
            15'd14341: log10_cal = 16'b0000010010010101;
            15'd14342: log10_cal = 16'b0000010010010101;
            15'd14343: log10_cal = 16'b0000010010010101;
            15'd14344: log10_cal = 16'b0000010010010101;
            15'd14345: log10_cal = 16'b0000010010010101;
            15'd14346: log10_cal = 16'b0000010010010101;
            15'd14347: log10_cal = 16'b0000010010010101;
            15'd14348: log10_cal = 16'b0000010010010110;
            15'd14349: log10_cal = 16'b0000010010010110;
            15'd14350: log10_cal = 16'b0000010010010110;
            15'd14351: log10_cal = 16'b0000010010010110;
            15'd14352: log10_cal = 16'b0000010010010110;
            15'd14353: log10_cal = 16'b0000010010010110;
            15'd14354: log10_cal = 16'b0000010010010110;
            15'd14355: log10_cal = 16'b0000010010010110;
            15'd14356: log10_cal = 16'b0000010010010110;
            15'd14357: log10_cal = 16'b0000010010010110;
            15'd14358: log10_cal = 16'b0000010010010110;
            15'd14359: log10_cal = 16'b0000010010010110;
            15'd14360: log10_cal = 16'b0000010010010110;
            15'd14361: log10_cal = 16'b0000010010010110;
            15'd14362: log10_cal = 16'b0000010010010110;
            15'd14363: log10_cal = 16'b0000010010010110;
            15'd14364: log10_cal = 16'b0000010010010110;
            15'd14365: log10_cal = 16'b0000010010010110;
            15'd14366: log10_cal = 16'b0000010010010110;
            15'd14367: log10_cal = 16'b0000010010010110;
            15'd14368: log10_cal = 16'b0000010010010110;
            15'd14369: log10_cal = 16'b0000010010010110;
            15'd14370: log10_cal = 16'b0000010010010110;
            15'd14371: log10_cal = 16'b0000010010010110;
            15'd14372: log10_cal = 16'b0000010010010110;
            15'd14373: log10_cal = 16'b0000010010010110;
            15'd14374: log10_cal = 16'b0000010010010110;
            15'd14375: log10_cal = 16'b0000010010010110;
            15'd14376: log10_cal = 16'b0000010010010110;
            15'd14377: log10_cal = 16'b0000010010010110;
            15'd14378: log10_cal = 16'b0000010010010110;
            15'd14379: log10_cal = 16'b0000010010010110;
            15'd14380: log10_cal = 16'b0000010010010110;
            15'd14381: log10_cal = 16'b0000010010010111;
            15'd14382: log10_cal = 16'b0000010010010111;
            15'd14383: log10_cal = 16'b0000010010010111;
            15'd14384: log10_cal = 16'b0000010010010111;
            15'd14385: log10_cal = 16'b0000010010010111;
            15'd14386: log10_cal = 16'b0000010010010111;
            15'd14387: log10_cal = 16'b0000010010010111;
            15'd14388: log10_cal = 16'b0000010010010111;
            15'd14389: log10_cal = 16'b0000010010010111;
            15'd14390: log10_cal = 16'b0000010010010111;
            15'd14391: log10_cal = 16'b0000010010010111;
            15'd14392: log10_cal = 16'b0000010010010111;
            15'd14393: log10_cal = 16'b0000010010010111;
            15'd14394: log10_cal = 16'b0000010010010111;
            15'd14395: log10_cal = 16'b0000010010010111;
            15'd14396: log10_cal = 16'b0000010010010111;
            15'd14397: log10_cal = 16'b0000010010010111;
            15'd14398: log10_cal = 16'b0000010010010111;
            15'd14399: log10_cal = 16'b0000010010010111;
            15'd14400: log10_cal = 16'b0000010010010111;
            15'd14401: log10_cal = 16'b0000010010010111;
            15'd14402: log10_cal = 16'b0000010010010111;
            15'd14403: log10_cal = 16'b0000010010010111;
            15'd14404: log10_cal = 16'b0000010010010111;
            15'd14405: log10_cal = 16'b0000010010010111;
            15'd14406: log10_cal = 16'b0000010010010111;
            15'd14407: log10_cal = 16'b0000010010010111;
            15'd14408: log10_cal = 16'b0000010010010111;
            15'd14409: log10_cal = 16'b0000010010010111;
            15'd14410: log10_cal = 16'b0000010010010111;
            15'd14411: log10_cal = 16'b0000010010010111;
            15'd14412: log10_cal = 16'b0000010010010111;
            15'd14413: log10_cal = 16'b0000010010011000;
            15'd14414: log10_cal = 16'b0000010010011000;
            15'd14415: log10_cal = 16'b0000010010011000;
            15'd14416: log10_cal = 16'b0000010010011000;
            15'd14417: log10_cal = 16'b0000010010011000;
            15'd14418: log10_cal = 16'b0000010010011000;
            15'd14419: log10_cal = 16'b0000010010011000;
            15'd14420: log10_cal = 16'b0000010010011000;
            15'd14421: log10_cal = 16'b0000010010011000;
            15'd14422: log10_cal = 16'b0000010010011000;
            15'd14423: log10_cal = 16'b0000010010011000;
            15'd14424: log10_cal = 16'b0000010010011000;
            15'd14425: log10_cal = 16'b0000010010011000;
            15'd14426: log10_cal = 16'b0000010010011000;
            15'd14427: log10_cal = 16'b0000010010011000;
            15'd14428: log10_cal = 16'b0000010010011000;
            15'd14429: log10_cal = 16'b0000010010011000;
            15'd14430: log10_cal = 16'b0000010010011000;
            15'd14431: log10_cal = 16'b0000010010011000;
            15'd14432: log10_cal = 16'b0000010010011000;
            15'd14433: log10_cal = 16'b0000010010011000;
            15'd14434: log10_cal = 16'b0000010010011000;
            15'd14435: log10_cal = 16'b0000010010011000;
            15'd14436: log10_cal = 16'b0000010010011000;
            15'd14437: log10_cal = 16'b0000010010011000;
            15'd14438: log10_cal = 16'b0000010010011000;
            15'd14439: log10_cal = 16'b0000010010011000;
            15'd14440: log10_cal = 16'b0000010010011000;
            15'd14441: log10_cal = 16'b0000010010011000;
            15'd14442: log10_cal = 16'b0000010010011000;
            15'd14443: log10_cal = 16'b0000010010011000;
            15'd14444: log10_cal = 16'b0000010010011000;
            15'd14445: log10_cal = 16'b0000010010011001;
            15'd14446: log10_cal = 16'b0000010010011001;
            15'd14447: log10_cal = 16'b0000010010011001;
            15'd14448: log10_cal = 16'b0000010010011001;
            15'd14449: log10_cal = 16'b0000010010011001;
            15'd14450: log10_cal = 16'b0000010010011001;
            15'd14451: log10_cal = 16'b0000010010011001;
            15'd14452: log10_cal = 16'b0000010010011001;
            15'd14453: log10_cal = 16'b0000010010011001;
            15'd14454: log10_cal = 16'b0000010010011001;
            15'd14455: log10_cal = 16'b0000010010011001;
            15'd14456: log10_cal = 16'b0000010010011001;
            15'd14457: log10_cal = 16'b0000010010011001;
            15'd14458: log10_cal = 16'b0000010010011001;
            15'd14459: log10_cal = 16'b0000010010011001;
            15'd14460: log10_cal = 16'b0000010010011001;
            15'd14461: log10_cal = 16'b0000010010011001;
            15'd14462: log10_cal = 16'b0000010010011001;
            15'd14463: log10_cal = 16'b0000010010011001;
            15'd14464: log10_cal = 16'b0000010010011001;
            15'd14465: log10_cal = 16'b0000010010011001;
            15'd14466: log10_cal = 16'b0000010010011001;
            15'd14467: log10_cal = 16'b0000010010011001;
            15'd14468: log10_cal = 16'b0000010010011001;
            15'd14469: log10_cal = 16'b0000010010011001;
            15'd14470: log10_cal = 16'b0000010010011001;
            15'd14471: log10_cal = 16'b0000010010011001;
            15'd14472: log10_cal = 16'b0000010010011001;
            15'd14473: log10_cal = 16'b0000010010011001;
            15'd14474: log10_cal = 16'b0000010010011001;
            15'd14475: log10_cal = 16'b0000010010011001;
            15'd14476: log10_cal = 16'b0000010010011001;
            15'd14477: log10_cal = 16'b0000010010011001;
            15'd14478: log10_cal = 16'b0000010010011010;
            15'd14479: log10_cal = 16'b0000010010011010;
            15'd14480: log10_cal = 16'b0000010010011010;
            15'd14481: log10_cal = 16'b0000010010011010;
            15'd14482: log10_cal = 16'b0000010010011010;
            15'd14483: log10_cal = 16'b0000010010011010;
            15'd14484: log10_cal = 16'b0000010010011010;
            15'd14485: log10_cal = 16'b0000010010011010;
            15'd14486: log10_cal = 16'b0000010010011010;
            15'd14487: log10_cal = 16'b0000010010011010;
            15'd14488: log10_cal = 16'b0000010010011010;
            15'd14489: log10_cal = 16'b0000010010011010;
            15'd14490: log10_cal = 16'b0000010010011010;
            15'd14491: log10_cal = 16'b0000010010011010;
            15'd14492: log10_cal = 16'b0000010010011010;
            15'd14493: log10_cal = 16'b0000010010011010;
            15'd14494: log10_cal = 16'b0000010010011010;
            15'd14495: log10_cal = 16'b0000010010011010;
            15'd14496: log10_cal = 16'b0000010010011010;
            15'd14497: log10_cal = 16'b0000010010011010;
            15'd14498: log10_cal = 16'b0000010010011010;
            15'd14499: log10_cal = 16'b0000010010011010;
            15'd14500: log10_cal = 16'b0000010010011010;
            15'd14501: log10_cal = 16'b0000010010011010;
            15'd14502: log10_cal = 16'b0000010010011010;
            15'd14503: log10_cal = 16'b0000010010011010;
            15'd14504: log10_cal = 16'b0000010010011010;
            15'd14505: log10_cal = 16'b0000010010011010;
            15'd14506: log10_cal = 16'b0000010010011010;
            15'd14507: log10_cal = 16'b0000010010011010;
            15'd14508: log10_cal = 16'b0000010010011010;
            15'd14509: log10_cal = 16'b0000010010011010;
            15'd14510: log10_cal = 16'b0000010010011011;
            15'd14511: log10_cal = 16'b0000010010011011;
            15'd14512: log10_cal = 16'b0000010010011011;
            15'd14513: log10_cal = 16'b0000010010011011;
            15'd14514: log10_cal = 16'b0000010010011011;
            15'd14515: log10_cal = 16'b0000010010011011;
            15'd14516: log10_cal = 16'b0000010010011011;
            15'd14517: log10_cal = 16'b0000010010011011;
            15'd14518: log10_cal = 16'b0000010010011011;
            15'd14519: log10_cal = 16'b0000010010011011;
            15'd14520: log10_cal = 16'b0000010010011011;
            15'd14521: log10_cal = 16'b0000010010011011;
            15'd14522: log10_cal = 16'b0000010010011011;
            15'd14523: log10_cal = 16'b0000010010011011;
            15'd14524: log10_cal = 16'b0000010010011011;
            15'd14525: log10_cal = 16'b0000010010011011;
            15'd14526: log10_cal = 16'b0000010010011011;
            15'd14527: log10_cal = 16'b0000010010011011;
            15'd14528: log10_cal = 16'b0000010010011011;
            15'd14529: log10_cal = 16'b0000010010011011;
            15'd14530: log10_cal = 16'b0000010010011011;
            15'd14531: log10_cal = 16'b0000010010011011;
            15'd14532: log10_cal = 16'b0000010010011011;
            15'd14533: log10_cal = 16'b0000010010011011;
            15'd14534: log10_cal = 16'b0000010010011011;
            15'd14535: log10_cal = 16'b0000010010011011;
            15'd14536: log10_cal = 16'b0000010010011011;
            15'd14537: log10_cal = 16'b0000010010011011;
            15'd14538: log10_cal = 16'b0000010010011011;
            15'd14539: log10_cal = 16'b0000010010011011;
            15'd14540: log10_cal = 16'b0000010010011011;
            15'd14541: log10_cal = 16'b0000010010011011;
            15'd14542: log10_cal = 16'b0000010010011011;
            15'd14543: log10_cal = 16'b0000010010011100;
            15'd14544: log10_cal = 16'b0000010010011100;
            15'd14545: log10_cal = 16'b0000010010011100;
            15'd14546: log10_cal = 16'b0000010010011100;
            15'd14547: log10_cal = 16'b0000010010011100;
            15'd14548: log10_cal = 16'b0000010010011100;
            15'd14549: log10_cal = 16'b0000010010011100;
            15'd14550: log10_cal = 16'b0000010010011100;
            15'd14551: log10_cal = 16'b0000010010011100;
            15'd14552: log10_cal = 16'b0000010010011100;
            15'd14553: log10_cal = 16'b0000010010011100;
            15'd14554: log10_cal = 16'b0000010010011100;
            15'd14555: log10_cal = 16'b0000010010011100;
            15'd14556: log10_cal = 16'b0000010010011100;
            15'd14557: log10_cal = 16'b0000010010011100;
            15'd14558: log10_cal = 16'b0000010010011100;
            15'd14559: log10_cal = 16'b0000010010011100;
            15'd14560: log10_cal = 16'b0000010010011100;
            15'd14561: log10_cal = 16'b0000010010011100;
            15'd14562: log10_cal = 16'b0000010010011100;
            15'd14563: log10_cal = 16'b0000010010011100;
            15'd14564: log10_cal = 16'b0000010010011100;
            15'd14565: log10_cal = 16'b0000010010011100;
            15'd14566: log10_cal = 16'b0000010010011100;
            15'd14567: log10_cal = 16'b0000010010011100;
            15'd14568: log10_cal = 16'b0000010010011100;
            15'd14569: log10_cal = 16'b0000010010011100;
            15'd14570: log10_cal = 16'b0000010010011100;
            15'd14571: log10_cal = 16'b0000010010011100;
            15'd14572: log10_cal = 16'b0000010010011100;
            15'd14573: log10_cal = 16'b0000010010011100;
            15'd14574: log10_cal = 16'b0000010010011100;
            15'd14575: log10_cal = 16'b0000010010011100;
            15'd14576: log10_cal = 16'b0000010010011101;
            15'd14577: log10_cal = 16'b0000010010011101;
            15'd14578: log10_cal = 16'b0000010010011101;
            15'd14579: log10_cal = 16'b0000010010011101;
            15'd14580: log10_cal = 16'b0000010010011101;
            15'd14581: log10_cal = 16'b0000010010011101;
            15'd14582: log10_cal = 16'b0000010010011101;
            15'd14583: log10_cal = 16'b0000010010011101;
            15'd14584: log10_cal = 16'b0000010010011101;
            15'd14585: log10_cal = 16'b0000010010011101;
            15'd14586: log10_cal = 16'b0000010010011101;
            15'd14587: log10_cal = 16'b0000010010011101;
            15'd14588: log10_cal = 16'b0000010010011101;
            15'd14589: log10_cal = 16'b0000010010011101;
            15'd14590: log10_cal = 16'b0000010010011101;
            15'd14591: log10_cal = 16'b0000010010011101;
            15'd14592: log10_cal = 16'b0000010010011101;
            15'd14593: log10_cal = 16'b0000010010011101;
            15'd14594: log10_cal = 16'b0000010010011101;
            15'd14595: log10_cal = 16'b0000010010011101;
            15'd14596: log10_cal = 16'b0000010010011101;
            15'd14597: log10_cal = 16'b0000010010011101;
            15'd14598: log10_cal = 16'b0000010010011101;
            15'd14599: log10_cal = 16'b0000010010011101;
            15'd14600: log10_cal = 16'b0000010010011101;
            15'd14601: log10_cal = 16'b0000010010011101;
            15'd14602: log10_cal = 16'b0000010010011101;
            15'd14603: log10_cal = 16'b0000010010011101;
            15'd14604: log10_cal = 16'b0000010010011101;
            15'd14605: log10_cal = 16'b0000010010011101;
            15'd14606: log10_cal = 16'b0000010010011101;
            15'd14607: log10_cal = 16'b0000010010011101;
            15'd14608: log10_cal = 16'b0000010010011101;
            15'd14609: log10_cal = 16'b0000010010011110;
            15'd14610: log10_cal = 16'b0000010010011110;
            15'd14611: log10_cal = 16'b0000010010011110;
            15'd14612: log10_cal = 16'b0000010010011110;
            15'd14613: log10_cal = 16'b0000010010011110;
            15'd14614: log10_cal = 16'b0000010010011110;
            15'd14615: log10_cal = 16'b0000010010011110;
            15'd14616: log10_cal = 16'b0000010010011110;
            15'd14617: log10_cal = 16'b0000010010011110;
            15'd14618: log10_cal = 16'b0000010010011110;
            15'd14619: log10_cal = 16'b0000010010011110;
            15'd14620: log10_cal = 16'b0000010010011110;
            15'd14621: log10_cal = 16'b0000010010011110;
            15'd14622: log10_cal = 16'b0000010010011110;
            15'd14623: log10_cal = 16'b0000010010011110;
            15'd14624: log10_cal = 16'b0000010010011110;
            15'd14625: log10_cal = 16'b0000010010011110;
            15'd14626: log10_cal = 16'b0000010010011110;
            15'd14627: log10_cal = 16'b0000010010011110;
            15'd14628: log10_cal = 16'b0000010010011110;
            15'd14629: log10_cal = 16'b0000010010011110;
            15'd14630: log10_cal = 16'b0000010010011110;
            15'd14631: log10_cal = 16'b0000010010011110;
            15'd14632: log10_cal = 16'b0000010010011110;
            15'd14633: log10_cal = 16'b0000010010011110;
            15'd14634: log10_cal = 16'b0000010010011110;
            15'd14635: log10_cal = 16'b0000010010011110;
            15'd14636: log10_cal = 16'b0000010010011110;
            15'd14637: log10_cal = 16'b0000010010011110;
            15'd14638: log10_cal = 16'b0000010010011110;
            15'd14639: log10_cal = 16'b0000010010011110;
            15'd14640: log10_cal = 16'b0000010010011110;
            15'd14641: log10_cal = 16'b0000010010011110;
            15'd14642: log10_cal = 16'b0000010010011111;
            15'd14643: log10_cal = 16'b0000010010011111;
            15'd14644: log10_cal = 16'b0000010010011111;
            15'd14645: log10_cal = 16'b0000010010011111;
            15'd14646: log10_cal = 16'b0000010010011111;
            15'd14647: log10_cal = 16'b0000010010011111;
            15'd14648: log10_cal = 16'b0000010010011111;
            15'd14649: log10_cal = 16'b0000010010011111;
            15'd14650: log10_cal = 16'b0000010010011111;
            15'd14651: log10_cal = 16'b0000010010011111;
            15'd14652: log10_cal = 16'b0000010010011111;
            15'd14653: log10_cal = 16'b0000010010011111;
            15'd14654: log10_cal = 16'b0000010010011111;
            15'd14655: log10_cal = 16'b0000010010011111;
            15'd14656: log10_cal = 16'b0000010010011111;
            15'd14657: log10_cal = 16'b0000010010011111;
            15'd14658: log10_cal = 16'b0000010010011111;
            15'd14659: log10_cal = 16'b0000010010011111;
            15'd14660: log10_cal = 16'b0000010010011111;
            15'd14661: log10_cal = 16'b0000010010011111;
            15'd14662: log10_cal = 16'b0000010010011111;
            15'd14663: log10_cal = 16'b0000010010011111;
            15'd14664: log10_cal = 16'b0000010010011111;
            15'd14665: log10_cal = 16'b0000010010011111;
            15'd14666: log10_cal = 16'b0000010010011111;
            15'd14667: log10_cal = 16'b0000010010011111;
            15'd14668: log10_cal = 16'b0000010010011111;
            15'd14669: log10_cal = 16'b0000010010011111;
            15'd14670: log10_cal = 16'b0000010010011111;
            15'd14671: log10_cal = 16'b0000010010011111;
            15'd14672: log10_cal = 16'b0000010010011111;
            15'd14673: log10_cal = 16'b0000010010011111;
            15'd14674: log10_cal = 16'b0000010010011111;
            15'd14675: log10_cal = 16'b0000010010100000;
            15'd14676: log10_cal = 16'b0000010010100000;
            15'd14677: log10_cal = 16'b0000010010100000;
            15'd14678: log10_cal = 16'b0000010010100000;
            15'd14679: log10_cal = 16'b0000010010100000;
            15'd14680: log10_cal = 16'b0000010010100000;
            15'd14681: log10_cal = 16'b0000010010100000;
            15'd14682: log10_cal = 16'b0000010010100000;
            15'd14683: log10_cal = 16'b0000010010100000;
            15'd14684: log10_cal = 16'b0000010010100000;
            15'd14685: log10_cal = 16'b0000010010100000;
            15'd14686: log10_cal = 16'b0000010010100000;
            15'd14687: log10_cal = 16'b0000010010100000;
            15'd14688: log10_cal = 16'b0000010010100000;
            15'd14689: log10_cal = 16'b0000010010100000;
            15'd14690: log10_cal = 16'b0000010010100000;
            15'd14691: log10_cal = 16'b0000010010100000;
            15'd14692: log10_cal = 16'b0000010010100000;
            15'd14693: log10_cal = 16'b0000010010100000;
            15'd14694: log10_cal = 16'b0000010010100000;
            15'd14695: log10_cal = 16'b0000010010100000;
            15'd14696: log10_cal = 16'b0000010010100000;
            15'd14697: log10_cal = 16'b0000010010100000;
            15'd14698: log10_cal = 16'b0000010010100000;
            15'd14699: log10_cal = 16'b0000010010100000;
            15'd14700: log10_cal = 16'b0000010010100000;
            15'd14701: log10_cal = 16'b0000010010100000;
            15'd14702: log10_cal = 16'b0000010010100000;
            15'd14703: log10_cal = 16'b0000010010100000;
            15'd14704: log10_cal = 16'b0000010010100000;
            15'd14705: log10_cal = 16'b0000010010100000;
            15'd14706: log10_cal = 16'b0000010010100000;
            15'd14707: log10_cal = 16'b0000010010100000;
            15'd14708: log10_cal = 16'b0000010010100001;
            15'd14709: log10_cal = 16'b0000010010100001;
            15'd14710: log10_cal = 16'b0000010010100001;
            15'd14711: log10_cal = 16'b0000010010100001;
            15'd14712: log10_cal = 16'b0000010010100001;
            15'd14713: log10_cal = 16'b0000010010100001;
            15'd14714: log10_cal = 16'b0000010010100001;
            15'd14715: log10_cal = 16'b0000010010100001;
            15'd14716: log10_cal = 16'b0000010010100001;
            15'd14717: log10_cal = 16'b0000010010100001;
            15'd14718: log10_cal = 16'b0000010010100001;
            15'd14719: log10_cal = 16'b0000010010100001;
            15'd14720: log10_cal = 16'b0000010010100001;
            15'd14721: log10_cal = 16'b0000010010100001;
            15'd14722: log10_cal = 16'b0000010010100001;
            15'd14723: log10_cal = 16'b0000010010100001;
            15'd14724: log10_cal = 16'b0000010010100001;
            15'd14725: log10_cal = 16'b0000010010100001;
            15'd14726: log10_cal = 16'b0000010010100001;
            15'd14727: log10_cal = 16'b0000010010100001;
            15'd14728: log10_cal = 16'b0000010010100001;
            15'd14729: log10_cal = 16'b0000010010100001;
            15'd14730: log10_cal = 16'b0000010010100001;
            15'd14731: log10_cal = 16'b0000010010100001;
            15'd14732: log10_cal = 16'b0000010010100001;
            15'd14733: log10_cal = 16'b0000010010100001;
            15'd14734: log10_cal = 16'b0000010010100001;
            15'd14735: log10_cal = 16'b0000010010100001;
            15'd14736: log10_cal = 16'b0000010010100001;
            15'd14737: log10_cal = 16'b0000010010100001;
            15'd14738: log10_cal = 16'b0000010010100001;
            15'd14739: log10_cal = 16'b0000010010100001;
            15'd14740: log10_cal = 16'b0000010010100001;
            15'd14741: log10_cal = 16'b0000010010100010;
            15'd14742: log10_cal = 16'b0000010010100010;
            15'd14743: log10_cal = 16'b0000010010100010;
            15'd14744: log10_cal = 16'b0000010010100010;
            15'd14745: log10_cal = 16'b0000010010100010;
            15'd14746: log10_cal = 16'b0000010010100010;
            15'd14747: log10_cal = 16'b0000010010100010;
            15'd14748: log10_cal = 16'b0000010010100010;
            15'd14749: log10_cal = 16'b0000010010100010;
            15'd14750: log10_cal = 16'b0000010010100010;
            15'd14751: log10_cal = 16'b0000010010100010;
            15'd14752: log10_cal = 16'b0000010010100010;
            15'd14753: log10_cal = 16'b0000010010100010;
            15'd14754: log10_cal = 16'b0000010010100010;
            15'd14755: log10_cal = 16'b0000010010100010;
            15'd14756: log10_cal = 16'b0000010010100010;
            15'd14757: log10_cal = 16'b0000010010100010;
            15'd14758: log10_cal = 16'b0000010010100010;
            15'd14759: log10_cal = 16'b0000010010100010;
            15'd14760: log10_cal = 16'b0000010010100010;
            15'd14761: log10_cal = 16'b0000010010100010;
            15'd14762: log10_cal = 16'b0000010010100010;
            15'd14763: log10_cal = 16'b0000010010100010;
            15'd14764: log10_cal = 16'b0000010010100010;
            15'd14765: log10_cal = 16'b0000010010100010;
            15'd14766: log10_cal = 16'b0000010010100010;
            15'd14767: log10_cal = 16'b0000010010100010;
            15'd14768: log10_cal = 16'b0000010010100010;
            15'd14769: log10_cal = 16'b0000010010100010;
            15'd14770: log10_cal = 16'b0000010010100010;
            15'd14771: log10_cal = 16'b0000010010100010;
            15'd14772: log10_cal = 16'b0000010010100010;
            15'd14773: log10_cal = 16'b0000010010100010;
            15'd14774: log10_cal = 16'b0000010010100011;
            15'd14775: log10_cal = 16'b0000010010100011;
            15'd14776: log10_cal = 16'b0000010010100011;
            15'd14777: log10_cal = 16'b0000010010100011;
            15'd14778: log10_cal = 16'b0000010010100011;
            15'd14779: log10_cal = 16'b0000010010100011;
            15'd14780: log10_cal = 16'b0000010010100011;
            15'd14781: log10_cal = 16'b0000010010100011;
            15'd14782: log10_cal = 16'b0000010010100011;
            15'd14783: log10_cal = 16'b0000010010100011;
            15'd14784: log10_cal = 16'b0000010010100011;
            15'd14785: log10_cal = 16'b0000010010100011;
            15'd14786: log10_cal = 16'b0000010010100011;
            15'd14787: log10_cal = 16'b0000010010100011;
            15'd14788: log10_cal = 16'b0000010010100011;
            15'd14789: log10_cal = 16'b0000010010100011;
            15'd14790: log10_cal = 16'b0000010010100011;
            15'd14791: log10_cal = 16'b0000010010100011;
            15'd14792: log10_cal = 16'b0000010010100011;
            15'd14793: log10_cal = 16'b0000010010100011;
            15'd14794: log10_cal = 16'b0000010010100011;
            15'd14795: log10_cal = 16'b0000010010100011;
            15'd14796: log10_cal = 16'b0000010010100011;
            15'd14797: log10_cal = 16'b0000010010100011;
            15'd14798: log10_cal = 16'b0000010010100011;
            15'd14799: log10_cal = 16'b0000010010100011;
            15'd14800: log10_cal = 16'b0000010010100011;
            15'd14801: log10_cal = 16'b0000010010100011;
            15'd14802: log10_cal = 16'b0000010010100011;
            15'd14803: log10_cal = 16'b0000010010100011;
            15'd14804: log10_cal = 16'b0000010010100011;
            15'd14805: log10_cal = 16'b0000010010100011;
            15'd14806: log10_cal = 16'b0000010010100011;
            15'd14807: log10_cal = 16'b0000010010100100;
            15'd14808: log10_cal = 16'b0000010010100100;
            15'd14809: log10_cal = 16'b0000010010100100;
            15'd14810: log10_cal = 16'b0000010010100100;
            15'd14811: log10_cal = 16'b0000010010100100;
            15'd14812: log10_cal = 16'b0000010010100100;
            15'd14813: log10_cal = 16'b0000010010100100;
            15'd14814: log10_cal = 16'b0000010010100100;
            15'd14815: log10_cal = 16'b0000010010100100;
            15'd14816: log10_cal = 16'b0000010010100100;
            15'd14817: log10_cal = 16'b0000010010100100;
            15'd14818: log10_cal = 16'b0000010010100100;
            15'd14819: log10_cal = 16'b0000010010100100;
            15'd14820: log10_cal = 16'b0000010010100100;
            15'd14821: log10_cal = 16'b0000010010100100;
            15'd14822: log10_cal = 16'b0000010010100100;
            15'd14823: log10_cal = 16'b0000010010100100;
            15'd14824: log10_cal = 16'b0000010010100100;
            15'd14825: log10_cal = 16'b0000010010100100;
            15'd14826: log10_cal = 16'b0000010010100100;
            15'd14827: log10_cal = 16'b0000010010100100;
            15'd14828: log10_cal = 16'b0000010010100100;
            15'd14829: log10_cal = 16'b0000010010100100;
            15'd14830: log10_cal = 16'b0000010010100100;
            15'd14831: log10_cal = 16'b0000010010100100;
            15'd14832: log10_cal = 16'b0000010010100100;
            15'd14833: log10_cal = 16'b0000010010100100;
            15'd14834: log10_cal = 16'b0000010010100100;
            15'd14835: log10_cal = 16'b0000010010100100;
            15'd14836: log10_cal = 16'b0000010010100100;
            15'd14837: log10_cal = 16'b0000010010100100;
            15'd14838: log10_cal = 16'b0000010010100100;
            15'd14839: log10_cal = 16'b0000010010100100;
            15'd14840: log10_cal = 16'b0000010010100101;
            15'd14841: log10_cal = 16'b0000010010100101;
            15'd14842: log10_cal = 16'b0000010010100101;
            15'd14843: log10_cal = 16'b0000010010100101;
            15'd14844: log10_cal = 16'b0000010010100101;
            15'd14845: log10_cal = 16'b0000010010100101;
            15'd14846: log10_cal = 16'b0000010010100101;
            15'd14847: log10_cal = 16'b0000010010100101;
            15'd14848: log10_cal = 16'b0000010010100101;
            15'd14849: log10_cal = 16'b0000010010100101;
            15'd14850: log10_cal = 16'b0000010010100101;
            15'd14851: log10_cal = 16'b0000010010100101;
            15'd14852: log10_cal = 16'b0000010010100101;
            15'd14853: log10_cal = 16'b0000010010100101;
            15'd14854: log10_cal = 16'b0000010010100101;
            15'd14855: log10_cal = 16'b0000010010100101;
            15'd14856: log10_cal = 16'b0000010010100101;
            15'd14857: log10_cal = 16'b0000010010100101;
            15'd14858: log10_cal = 16'b0000010010100101;
            15'd14859: log10_cal = 16'b0000010010100101;
            15'd14860: log10_cal = 16'b0000010010100101;
            15'd14861: log10_cal = 16'b0000010010100101;
            15'd14862: log10_cal = 16'b0000010010100101;
            15'd14863: log10_cal = 16'b0000010010100101;
            15'd14864: log10_cal = 16'b0000010010100101;
            15'd14865: log10_cal = 16'b0000010010100101;
            15'd14866: log10_cal = 16'b0000010010100101;
            15'd14867: log10_cal = 16'b0000010010100101;
            15'd14868: log10_cal = 16'b0000010010100101;
            15'd14869: log10_cal = 16'b0000010010100101;
            15'd14870: log10_cal = 16'b0000010010100101;
            15'd14871: log10_cal = 16'b0000010010100101;
            15'd14872: log10_cal = 16'b0000010010100101;
            15'd14873: log10_cal = 16'b0000010010100101;
            15'd14874: log10_cal = 16'b0000010010100110;
            15'd14875: log10_cal = 16'b0000010010100110;
            15'd14876: log10_cal = 16'b0000010010100110;
            15'd14877: log10_cal = 16'b0000010010100110;
            15'd14878: log10_cal = 16'b0000010010100110;
            15'd14879: log10_cal = 16'b0000010010100110;
            15'd14880: log10_cal = 16'b0000010010100110;
            15'd14881: log10_cal = 16'b0000010010100110;
            15'd14882: log10_cal = 16'b0000010010100110;
            15'd14883: log10_cal = 16'b0000010010100110;
            15'd14884: log10_cal = 16'b0000010010100110;
            15'd14885: log10_cal = 16'b0000010010100110;
            15'd14886: log10_cal = 16'b0000010010100110;
            15'd14887: log10_cal = 16'b0000010010100110;
            15'd14888: log10_cal = 16'b0000010010100110;
            15'd14889: log10_cal = 16'b0000010010100110;
            15'd14890: log10_cal = 16'b0000010010100110;
            15'd14891: log10_cal = 16'b0000010010100110;
            15'd14892: log10_cal = 16'b0000010010100110;
            15'd14893: log10_cal = 16'b0000010010100110;
            15'd14894: log10_cal = 16'b0000010010100110;
            15'd14895: log10_cal = 16'b0000010010100110;
            15'd14896: log10_cal = 16'b0000010010100110;
            15'd14897: log10_cal = 16'b0000010010100110;
            15'd14898: log10_cal = 16'b0000010010100110;
            15'd14899: log10_cal = 16'b0000010010100110;
            15'd14900: log10_cal = 16'b0000010010100110;
            15'd14901: log10_cal = 16'b0000010010100110;
            15'd14902: log10_cal = 16'b0000010010100110;
            15'd14903: log10_cal = 16'b0000010010100110;
            15'd14904: log10_cal = 16'b0000010010100110;
            15'd14905: log10_cal = 16'b0000010010100110;
            15'd14906: log10_cal = 16'b0000010010100110;
            15'd14907: log10_cal = 16'b0000010010100111;
            15'd14908: log10_cal = 16'b0000010010100111;
            15'd14909: log10_cal = 16'b0000010010100111;
            15'd14910: log10_cal = 16'b0000010010100111;
            15'd14911: log10_cal = 16'b0000010010100111;
            15'd14912: log10_cal = 16'b0000010010100111;
            15'd14913: log10_cal = 16'b0000010010100111;
            15'd14914: log10_cal = 16'b0000010010100111;
            15'd14915: log10_cal = 16'b0000010010100111;
            15'd14916: log10_cal = 16'b0000010010100111;
            15'd14917: log10_cal = 16'b0000010010100111;
            15'd14918: log10_cal = 16'b0000010010100111;
            15'd14919: log10_cal = 16'b0000010010100111;
            15'd14920: log10_cal = 16'b0000010010100111;
            15'd14921: log10_cal = 16'b0000010010100111;
            15'd14922: log10_cal = 16'b0000010010100111;
            15'd14923: log10_cal = 16'b0000010010100111;
            15'd14924: log10_cal = 16'b0000010010100111;
            15'd14925: log10_cal = 16'b0000010010100111;
            15'd14926: log10_cal = 16'b0000010010100111;
            15'd14927: log10_cal = 16'b0000010010100111;
            15'd14928: log10_cal = 16'b0000010010100111;
            15'd14929: log10_cal = 16'b0000010010100111;
            15'd14930: log10_cal = 16'b0000010010100111;
            15'd14931: log10_cal = 16'b0000010010100111;
            15'd14932: log10_cal = 16'b0000010010100111;
            15'd14933: log10_cal = 16'b0000010010100111;
            15'd14934: log10_cal = 16'b0000010010100111;
            15'd14935: log10_cal = 16'b0000010010100111;
            15'd14936: log10_cal = 16'b0000010010100111;
            15'd14937: log10_cal = 16'b0000010010100111;
            15'd14938: log10_cal = 16'b0000010010100111;
            15'd14939: log10_cal = 16'b0000010010100111;
            15'd14940: log10_cal = 16'b0000010010100111;
            15'd14941: log10_cal = 16'b0000010010101000;
            15'd14942: log10_cal = 16'b0000010010101000;
            15'd14943: log10_cal = 16'b0000010010101000;
            15'd14944: log10_cal = 16'b0000010010101000;
            15'd14945: log10_cal = 16'b0000010010101000;
            15'd14946: log10_cal = 16'b0000010010101000;
            15'd14947: log10_cal = 16'b0000010010101000;
            15'd14948: log10_cal = 16'b0000010010101000;
            15'd14949: log10_cal = 16'b0000010010101000;
            15'd14950: log10_cal = 16'b0000010010101000;
            15'd14951: log10_cal = 16'b0000010010101000;
            15'd14952: log10_cal = 16'b0000010010101000;
            15'd14953: log10_cal = 16'b0000010010101000;
            15'd14954: log10_cal = 16'b0000010010101000;
            15'd14955: log10_cal = 16'b0000010010101000;
            15'd14956: log10_cal = 16'b0000010010101000;
            15'd14957: log10_cal = 16'b0000010010101000;
            15'd14958: log10_cal = 16'b0000010010101000;
            15'd14959: log10_cal = 16'b0000010010101000;
            15'd14960: log10_cal = 16'b0000010010101000;
            15'd14961: log10_cal = 16'b0000010010101000;
            15'd14962: log10_cal = 16'b0000010010101000;
            15'd14963: log10_cal = 16'b0000010010101000;
            15'd14964: log10_cal = 16'b0000010010101000;
            15'd14965: log10_cal = 16'b0000010010101000;
            15'd14966: log10_cal = 16'b0000010010101000;
            15'd14967: log10_cal = 16'b0000010010101000;
            15'd14968: log10_cal = 16'b0000010010101000;
            15'd14969: log10_cal = 16'b0000010010101000;
            15'd14970: log10_cal = 16'b0000010010101000;
            15'd14971: log10_cal = 16'b0000010010101000;
            15'd14972: log10_cal = 16'b0000010010101000;
            15'd14973: log10_cal = 16'b0000010010101000;
            15'd14974: log10_cal = 16'b0000010010101000;
            15'd14975: log10_cal = 16'b0000010010101001;
            15'd14976: log10_cal = 16'b0000010010101001;
            15'd14977: log10_cal = 16'b0000010010101001;
            15'd14978: log10_cal = 16'b0000010010101001;
            15'd14979: log10_cal = 16'b0000010010101001;
            15'd14980: log10_cal = 16'b0000010010101001;
            15'd14981: log10_cal = 16'b0000010010101001;
            15'd14982: log10_cal = 16'b0000010010101001;
            15'd14983: log10_cal = 16'b0000010010101001;
            15'd14984: log10_cal = 16'b0000010010101001;
            15'd14985: log10_cal = 16'b0000010010101001;
            15'd14986: log10_cal = 16'b0000010010101001;
            15'd14987: log10_cal = 16'b0000010010101001;
            15'd14988: log10_cal = 16'b0000010010101001;
            15'd14989: log10_cal = 16'b0000010010101001;
            15'd14990: log10_cal = 16'b0000010010101001;
            15'd14991: log10_cal = 16'b0000010010101001;
            15'd14992: log10_cal = 16'b0000010010101001;
            15'd14993: log10_cal = 16'b0000010010101001;
            15'd14994: log10_cal = 16'b0000010010101001;
            15'd14995: log10_cal = 16'b0000010010101001;
            15'd14996: log10_cal = 16'b0000010010101001;
            15'd14997: log10_cal = 16'b0000010010101001;
            15'd14998: log10_cal = 16'b0000010010101001;
            15'd14999: log10_cal = 16'b0000010010101001;
            15'd15000: log10_cal = 16'b0000010010101001;
            15'd15001: log10_cal = 16'b0000010010101001;
            15'd15002: log10_cal = 16'b0000010010101001;
            15'd15003: log10_cal = 16'b0000010010101001;
            15'd15004: log10_cal = 16'b0000010010101001;
            15'd15005: log10_cal = 16'b0000010010101001;
            15'd15006: log10_cal = 16'b0000010010101001;
            15'd15007: log10_cal = 16'b0000010010101001;
            15'd15008: log10_cal = 16'b0000010010101010;
            15'd15009: log10_cal = 16'b0000010010101010;
            15'd15010: log10_cal = 16'b0000010010101010;
            15'd15011: log10_cal = 16'b0000010010101010;
            15'd15012: log10_cal = 16'b0000010010101010;
            15'd15013: log10_cal = 16'b0000010010101010;
            15'd15014: log10_cal = 16'b0000010010101010;
            15'd15015: log10_cal = 16'b0000010010101010;
            15'd15016: log10_cal = 16'b0000010010101010;
            15'd15017: log10_cal = 16'b0000010010101010;
            15'd15018: log10_cal = 16'b0000010010101010;
            15'd15019: log10_cal = 16'b0000010010101010;
            15'd15020: log10_cal = 16'b0000010010101010;
            15'd15021: log10_cal = 16'b0000010010101010;
            15'd15022: log10_cal = 16'b0000010010101010;
            15'd15023: log10_cal = 16'b0000010010101010;
            15'd15024: log10_cal = 16'b0000010010101010;
            15'd15025: log10_cal = 16'b0000010010101010;
            15'd15026: log10_cal = 16'b0000010010101010;
            15'd15027: log10_cal = 16'b0000010010101010;
            15'd15028: log10_cal = 16'b0000010010101010;
            15'd15029: log10_cal = 16'b0000010010101010;
            15'd15030: log10_cal = 16'b0000010010101010;
            15'd15031: log10_cal = 16'b0000010010101010;
            15'd15032: log10_cal = 16'b0000010010101010;
            15'd15033: log10_cal = 16'b0000010010101010;
            15'd15034: log10_cal = 16'b0000010010101010;
            15'd15035: log10_cal = 16'b0000010010101010;
            15'd15036: log10_cal = 16'b0000010010101010;
            15'd15037: log10_cal = 16'b0000010010101010;
            15'd15038: log10_cal = 16'b0000010010101010;
            15'd15039: log10_cal = 16'b0000010010101010;
            15'd15040: log10_cal = 16'b0000010010101010;
            15'd15041: log10_cal = 16'b0000010010101010;
            15'd15042: log10_cal = 16'b0000010010101011;
            15'd15043: log10_cal = 16'b0000010010101011;
            15'd15044: log10_cal = 16'b0000010010101011;
            15'd15045: log10_cal = 16'b0000010010101011;
            15'd15046: log10_cal = 16'b0000010010101011;
            15'd15047: log10_cal = 16'b0000010010101011;
            15'd15048: log10_cal = 16'b0000010010101011;
            15'd15049: log10_cal = 16'b0000010010101011;
            15'd15050: log10_cal = 16'b0000010010101011;
            15'd15051: log10_cal = 16'b0000010010101011;
            15'd15052: log10_cal = 16'b0000010010101011;
            15'd15053: log10_cal = 16'b0000010010101011;
            15'd15054: log10_cal = 16'b0000010010101011;
            15'd15055: log10_cal = 16'b0000010010101011;
            15'd15056: log10_cal = 16'b0000010010101011;
            15'd15057: log10_cal = 16'b0000010010101011;
            15'd15058: log10_cal = 16'b0000010010101011;
            15'd15059: log10_cal = 16'b0000010010101011;
            15'd15060: log10_cal = 16'b0000010010101011;
            15'd15061: log10_cal = 16'b0000010010101011;
            15'd15062: log10_cal = 16'b0000010010101011;
            15'd15063: log10_cal = 16'b0000010010101011;
            15'd15064: log10_cal = 16'b0000010010101011;
            15'd15065: log10_cal = 16'b0000010010101011;
            15'd15066: log10_cal = 16'b0000010010101011;
            15'd15067: log10_cal = 16'b0000010010101011;
            15'd15068: log10_cal = 16'b0000010010101011;
            15'd15069: log10_cal = 16'b0000010010101011;
            15'd15070: log10_cal = 16'b0000010010101011;
            15'd15071: log10_cal = 16'b0000010010101011;
            15'd15072: log10_cal = 16'b0000010010101011;
            15'd15073: log10_cal = 16'b0000010010101011;
            15'd15074: log10_cal = 16'b0000010010101011;
            15'd15075: log10_cal = 16'b0000010010101011;
            15'd15076: log10_cal = 16'b0000010010101100;
            15'd15077: log10_cal = 16'b0000010010101100;
            15'd15078: log10_cal = 16'b0000010010101100;
            15'd15079: log10_cal = 16'b0000010010101100;
            15'd15080: log10_cal = 16'b0000010010101100;
            15'd15081: log10_cal = 16'b0000010010101100;
            15'd15082: log10_cal = 16'b0000010010101100;
            15'd15083: log10_cal = 16'b0000010010101100;
            15'd15084: log10_cal = 16'b0000010010101100;
            15'd15085: log10_cal = 16'b0000010010101100;
            15'd15086: log10_cal = 16'b0000010010101100;
            15'd15087: log10_cal = 16'b0000010010101100;
            15'd15088: log10_cal = 16'b0000010010101100;
            15'd15089: log10_cal = 16'b0000010010101100;
            15'd15090: log10_cal = 16'b0000010010101100;
            15'd15091: log10_cal = 16'b0000010010101100;
            15'd15092: log10_cal = 16'b0000010010101100;
            15'd15093: log10_cal = 16'b0000010010101100;
            15'd15094: log10_cal = 16'b0000010010101100;
            15'd15095: log10_cal = 16'b0000010010101100;
            15'd15096: log10_cal = 16'b0000010010101100;
            15'd15097: log10_cal = 16'b0000010010101100;
            15'd15098: log10_cal = 16'b0000010010101100;
            15'd15099: log10_cal = 16'b0000010010101100;
            15'd15100: log10_cal = 16'b0000010010101100;
            15'd15101: log10_cal = 16'b0000010010101100;
            15'd15102: log10_cal = 16'b0000010010101100;
            15'd15103: log10_cal = 16'b0000010010101100;
            15'd15104: log10_cal = 16'b0000010010101100;
            15'd15105: log10_cal = 16'b0000010010101100;
            15'd15106: log10_cal = 16'b0000010010101100;
            15'd15107: log10_cal = 16'b0000010010101100;
            15'd15108: log10_cal = 16'b0000010010101100;
            15'd15109: log10_cal = 16'b0000010010101100;
            15'd15110: log10_cal = 16'b0000010010101101;
            15'd15111: log10_cal = 16'b0000010010101101;
            15'd15112: log10_cal = 16'b0000010010101101;
            15'd15113: log10_cal = 16'b0000010010101101;
            15'd15114: log10_cal = 16'b0000010010101101;
            15'd15115: log10_cal = 16'b0000010010101101;
            15'd15116: log10_cal = 16'b0000010010101101;
            15'd15117: log10_cal = 16'b0000010010101101;
            15'd15118: log10_cal = 16'b0000010010101101;
            15'd15119: log10_cal = 16'b0000010010101101;
            15'd15120: log10_cal = 16'b0000010010101101;
            15'd15121: log10_cal = 16'b0000010010101101;
            15'd15122: log10_cal = 16'b0000010010101101;
            15'd15123: log10_cal = 16'b0000010010101101;
            15'd15124: log10_cal = 16'b0000010010101101;
            15'd15125: log10_cal = 16'b0000010010101101;
            15'd15126: log10_cal = 16'b0000010010101101;
            15'd15127: log10_cal = 16'b0000010010101101;
            15'd15128: log10_cal = 16'b0000010010101101;
            15'd15129: log10_cal = 16'b0000010010101101;
            15'd15130: log10_cal = 16'b0000010010101101;
            15'd15131: log10_cal = 16'b0000010010101101;
            15'd15132: log10_cal = 16'b0000010010101101;
            15'd15133: log10_cal = 16'b0000010010101101;
            15'd15134: log10_cal = 16'b0000010010101101;
            15'd15135: log10_cal = 16'b0000010010101101;
            15'd15136: log10_cal = 16'b0000010010101101;
            15'd15137: log10_cal = 16'b0000010010101101;
            15'd15138: log10_cal = 16'b0000010010101101;
            15'd15139: log10_cal = 16'b0000010010101101;
            15'd15140: log10_cal = 16'b0000010010101101;
            15'd15141: log10_cal = 16'b0000010010101101;
            15'd15142: log10_cal = 16'b0000010010101101;
            15'd15143: log10_cal = 16'b0000010010101101;
            15'd15144: log10_cal = 16'b0000010010101110;
            15'd15145: log10_cal = 16'b0000010010101110;
            15'd15146: log10_cal = 16'b0000010010101110;
            15'd15147: log10_cal = 16'b0000010010101110;
            15'd15148: log10_cal = 16'b0000010010101110;
            15'd15149: log10_cal = 16'b0000010010101110;
            15'd15150: log10_cal = 16'b0000010010101110;
            15'd15151: log10_cal = 16'b0000010010101110;
            15'd15152: log10_cal = 16'b0000010010101110;
            15'd15153: log10_cal = 16'b0000010010101110;
            15'd15154: log10_cal = 16'b0000010010101110;
            15'd15155: log10_cal = 16'b0000010010101110;
            15'd15156: log10_cal = 16'b0000010010101110;
            15'd15157: log10_cal = 16'b0000010010101110;
            15'd15158: log10_cal = 16'b0000010010101110;
            15'd15159: log10_cal = 16'b0000010010101110;
            15'd15160: log10_cal = 16'b0000010010101110;
            15'd15161: log10_cal = 16'b0000010010101110;
            15'd15162: log10_cal = 16'b0000010010101110;
            15'd15163: log10_cal = 16'b0000010010101110;
            15'd15164: log10_cal = 16'b0000010010101110;
            15'd15165: log10_cal = 16'b0000010010101110;
            15'd15166: log10_cal = 16'b0000010010101110;
            15'd15167: log10_cal = 16'b0000010010101110;
            15'd15168: log10_cal = 16'b0000010010101110;
            15'd15169: log10_cal = 16'b0000010010101110;
            15'd15170: log10_cal = 16'b0000010010101110;
            15'd15171: log10_cal = 16'b0000010010101110;
            15'd15172: log10_cal = 16'b0000010010101110;
            15'd15173: log10_cal = 16'b0000010010101110;
            15'd15174: log10_cal = 16'b0000010010101110;
            15'd15175: log10_cal = 16'b0000010010101110;
            15'd15176: log10_cal = 16'b0000010010101110;
            15'd15177: log10_cal = 16'b0000010010101110;
            15'd15178: log10_cal = 16'b0000010010101111;
            15'd15179: log10_cal = 16'b0000010010101111;
            15'd15180: log10_cal = 16'b0000010010101111;
            15'd15181: log10_cal = 16'b0000010010101111;
            15'd15182: log10_cal = 16'b0000010010101111;
            15'd15183: log10_cal = 16'b0000010010101111;
            15'd15184: log10_cal = 16'b0000010010101111;
            15'd15185: log10_cal = 16'b0000010010101111;
            15'd15186: log10_cal = 16'b0000010010101111;
            15'd15187: log10_cal = 16'b0000010010101111;
            15'd15188: log10_cal = 16'b0000010010101111;
            15'd15189: log10_cal = 16'b0000010010101111;
            15'd15190: log10_cal = 16'b0000010010101111;
            15'd15191: log10_cal = 16'b0000010010101111;
            15'd15192: log10_cal = 16'b0000010010101111;
            15'd15193: log10_cal = 16'b0000010010101111;
            15'd15194: log10_cal = 16'b0000010010101111;
            15'd15195: log10_cal = 16'b0000010010101111;
            15'd15196: log10_cal = 16'b0000010010101111;
            15'd15197: log10_cal = 16'b0000010010101111;
            15'd15198: log10_cal = 16'b0000010010101111;
            15'd15199: log10_cal = 16'b0000010010101111;
            15'd15200: log10_cal = 16'b0000010010101111;
            15'd15201: log10_cal = 16'b0000010010101111;
            15'd15202: log10_cal = 16'b0000010010101111;
            15'd15203: log10_cal = 16'b0000010010101111;
            15'd15204: log10_cal = 16'b0000010010101111;
            15'd15205: log10_cal = 16'b0000010010101111;
            15'd15206: log10_cal = 16'b0000010010101111;
            15'd15207: log10_cal = 16'b0000010010101111;
            15'd15208: log10_cal = 16'b0000010010101111;
            15'd15209: log10_cal = 16'b0000010010101111;
            15'd15210: log10_cal = 16'b0000010010101111;
            15'd15211: log10_cal = 16'b0000010010101111;
            15'd15212: log10_cal = 16'b0000010010110000;
            15'd15213: log10_cal = 16'b0000010010110000;
            15'd15214: log10_cal = 16'b0000010010110000;
            15'd15215: log10_cal = 16'b0000010010110000;
            15'd15216: log10_cal = 16'b0000010010110000;
            15'd15217: log10_cal = 16'b0000010010110000;
            15'd15218: log10_cal = 16'b0000010010110000;
            15'd15219: log10_cal = 16'b0000010010110000;
            15'd15220: log10_cal = 16'b0000010010110000;
            15'd15221: log10_cal = 16'b0000010010110000;
            15'd15222: log10_cal = 16'b0000010010110000;
            15'd15223: log10_cal = 16'b0000010010110000;
            15'd15224: log10_cal = 16'b0000010010110000;
            15'd15225: log10_cal = 16'b0000010010110000;
            15'd15226: log10_cal = 16'b0000010010110000;
            15'd15227: log10_cal = 16'b0000010010110000;
            15'd15228: log10_cal = 16'b0000010010110000;
            15'd15229: log10_cal = 16'b0000010010110000;
            15'd15230: log10_cal = 16'b0000010010110000;
            15'd15231: log10_cal = 16'b0000010010110000;
            15'd15232: log10_cal = 16'b0000010010110000;
            15'd15233: log10_cal = 16'b0000010010110000;
            15'd15234: log10_cal = 16'b0000010010110000;
            15'd15235: log10_cal = 16'b0000010010110000;
            15'd15236: log10_cal = 16'b0000010010110000;
            15'd15237: log10_cal = 16'b0000010010110000;
            15'd15238: log10_cal = 16'b0000010010110000;
            15'd15239: log10_cal = 16'b0000010010110000;
            15'd15240: log10_cal = 16'b0000010010110000;
            15'd15241: log10_cal = 16'b0000010010110000;
            15'd15242: log10_cal = 16'b0000010010110000;
            15'd15243: log10_cal = 16'b0000010010110000;
            15'd15244: log10_cal = 16'b0000010010110000;
            15'd15245: log10_cal = 16'b0000010010110000;
            15'd15246: log10_cal = 16'b0000010010110001;
            15'd15247: log10_cal = 16'b0000010010110001;
            15'd15248: log10_cal = 16'b0000010010110001;
            15'd15249: log10_cal = 16'b0000010010110001;
            15'd15250: log10_cal = 16'b0000010010110001;
            15'd15251: log10_cal = 16'b0000010010110001;
            15'd15252: log10_cal = 16'b0000010010110001;
            15'd15253: log10_cal = 16'b0000010010110001;
            15'd15254: log10_cal = 16'b0000010010110001;
            15'd15255: log10_cal = 16'b0000010010110001;
            15'd15256: log10_cal = 16'b0000010010110001;
            15'd15257: log10_cal = 16'b0000010010110001;
            15'd15258: log10_cal = 16'b0000010010110001;
            15'd15259: log10_cal = 16'b0000010010110001;
            15'd15260: log10_cal = 16'b0000010010110001;
            15'd15261: log10_cal = 16'b0000010010110001;
            15'd15262: log10_cal = 16'b0000010010110001;
            15'd15263: log10_cal = 16'b0000010010110001;
            15'd15264: log10_cal = 16'b0000010010110001;
            15'd15265: log10_cal = 16'b0000010010110001;
            15'd15266: log10_cal = 16'b0000010010110001;
            15'd15267: log10_cal = 16'b0000010010110001;
            15'd15268: log10_cal = 16'b0000010010110001;
            15'd15269: log10_cal = 16'b0000010010110001;
            15'd15270: log10_cal = 16'b0000010010110001;
            15'd15271: log10_cal = 16'b0000010010110001;
            15'd15272: log10_cal = 16'b0000010010110001;
            15'd15273: log10_cal = 16'b0000010010110001;
            15'd15274: log10_cal = 16'b0000010010110001;
            15'd15275: log10_cal = 16'b0000010010110001;
            15'd15276: log10_cal = 16'b0000010010110001;
            15'd15277: log10_cal = 16'b0000010010110001;
            15'd15278: log10_cal = 16'b0000010010110001;
            15'd15279: log10_cal = 16'b0000010010110001;
            15'd15280: log10_cal = 16'b0000010010110001;
            15'd15281: log10_cal = 16'b0000010010110010;
            15'd15282: log10_cal = 16'b0000010010110010;
            15'd15283: log10_cal = 16'b0000010010110010;
            15'd15284: log10_cal = 16'b0000010010110010;
            15'd15285: log10_cal = 16'b0000010010110010;
            15'd15286: log10_cal = 16'b0000010010110010;
            15'd15287: log10_cal = 16'b0000010010110010;
            15'd15288: log10_cal = 16'b0000010010110010;
            15'd15289: log10_cal = 16'b0000010010110010;
            15'd15290: log10_cal = 16'b0000010010110010;
            15'd15291: log10_cal = 16'b0000010010110010;
            15'd15292: log10_cal = 16'b0000010010110010;
            15'd15293: log10_cal = 16'b0000010010110010;
            15'd15294: log10_cal = 16'b0000010010110010;
            15'd15295: log10_cal = 16'b0000010010110010;
            15'd15296: log10_cal = 16'b0000010010110010;
            15'd15297: log10_cal = 16'b0000010010110010;
            15'd15298: log10_cal = 16'b0000010010110010;
            15'd15299: log10_cal = 16'b0000010010110010;
            15'd15300: log10_cal = 16'b0000010010110010;
            15'd15301: log10_cal = 16'b0000010010110010;
            15'd15302: log10_cal = 16'b0000010010110010;
            15'd15303: log10_cal = 16'b0000010010110010;
            15'd15304: log10_cal = 16'b0000010010110010;
            15'd15305: log10_cal = 16'b0000010010110010;
            15'd15306: log10_cal = 16'b0000010010110010;
            15'd15307: log10_cal = 16'b0000010010110010;
            15'd15308: log10_cal = 16'b0000010010110010;
            15'd15309: log10_cal = 16'b0000010010110010;
            15'd15310: log10_cal = 16'b0000010010110010;
            15'd15311: log10_cal = 16'b0000010010110010;
            15'd15312: log10_cal = 16'b0000010010110010;
            15'd15313: log10_cal = 16'b0000010010110010;
            15'd15314: log10_cal = 16'b0000010010110010;
            15'd15315: log10_cal = 16'b0000010010110011;
            15'd15316: log10_cal = 16'b0000010010110011;
            15'd15317: log10_cal = 16'b0000010010110011;
            15'd15318: log10_cal = 16'b0000010010110011;
            15'd15319: log10_cal = 16'b0000010010110011;
            15'd15320: log10_cal = 16'b0000010010110011;
            15'd15321: log10_cal = 16'b0000010010110011;
            15'd15322: log10_cal = 16'b0000010010110011;
            15'd15323: log10_cal = 16'b0000010010110011;
            15'd15324: log10_cal = 16'b0000010010110011;
            15'd15325: log10_cal = 16'b0000010010110011;
            15'd15326: log10_cal = 16'b0000010010110011;
            15'd15327: log10_cal = 16'b0000010010110011;
            15'd15328: log10_cal = 16'b0000010010110011;
            15'd15329: log10_cal = 16'b0000010010110011;
            15'd15330: log10_cal = 16'b0000010010110011;
            15'd15331: log10_cal = 16'b0000010010110011;
            15'd15332: log10_cal = 16'b0000010010110011;
            15'd15333: log10_cal = 16'b0000010010110011;
            15'd15334: log10_cal = 16'b0000010010110011;
            15'd15335: log10_cal = 16'b0000010010110011;
            15'd15336: log10_cal = 16'b0000010010110011;
            15'd15337: log10_cal = 16'b0000010010110011;
            15'd15338: log10_cal = 16'b0000010010110011;
            15'd15339: log10_cal = 16'b0000010010110011;
            15'd15340: log10_cal = 16'b0000010010110011;
            15'd15341: log10_cal = 16'b0000010010110011;
            15'd15342: log10_cal = 16'b0000010010110011;
            15'd15343: log10_cal = 16'b0000010010110011;
            15'd15344: log10_cal = 16'b0000010010110011;
            15'd15345: log10_cal = 16'b0000010010110011;
            15'd15346: log10_cal = 16'b0000010010110011;
            15'd15347: log10_cal = 16'b0000010010110011;
            15'd15348: log10_cal = 16'b0000010010110011;
            15'd15349: log10_cal = 16'b0000010010110011;
            15'd15350: log10_cal = 16'b0000010010110100;
            15'd15351: log10_cal = 16'b0000010010110100;
            15'd15352: log10_cal = 16'b0000010010110100;
            15'd15353: log10_cal = 16'b0000010010110100;
            15'd15354: log10_cal = 16'b0000010010110100;
            15'd15355: log10_cal = 16'b0000010010110100;
            15'd15356: log10_cal = 16'b0000010010110100;
            15'd15357: log10_cal = 16'b0000010010110100;
            15'd15358: log10_cal = 16'b0000010010110100;
            15'd15359: log10_cal = 16'b0000010010110100;
            15'd15360: log10_cal = 16'b0000010010110100;
            15'd15361: log10_cal = 16'b0000010010110100;
            15'd15362: log10_cal = 16'b0000010010110100;
            15'd15363: log10_cal = 16'b0000010010110100;
            15'd15364: log10_cal = 16'b0000010010110100;
            15'd15365: log10_cal = 16'b0000010010110100;
            15'd15366: log10_cal = 16'b0000010010110100;
            15'd15367: log10_cal = 16'b0000010010110100;
            15'd15368: log10_cal = 16'b0000010010110100;
            15'd15369: log10_cal = 16'b0000010010110100;
            15'd15370: log10_cal = 16'b0000010010110100;
            15'd15371: log10_cal = 16'b0000010010110100;
            15'd15372: log10_cal = 16'b0000010010110100;
            15'd15373: log10_cal = 16'b0000010010110100;
            15'd15374: log10_cal = 16'b0000010010110100;
            15'd15375: log10_cal = 16'b0000010010110100;
            15'd15376: log10_cal = 16'b0000010010110100;
            15'd15377: log10_cal = 16'b0000010010110100;
            15'd15378: log10_cal = 16'b0000010010110100;
            15'd15379: log10_cal = 16'b0000010010110100;
            15'd15380: log10_cal = 16'b0000010010110100;
            15'd15381: log10_cal = 16'b0000010010110100;
            15'd15382: log10_cal = 16'b0000010010110100;
            15'd15383: log10_cal = 16'b0000010010110100;
            15'd15384: log10_cal = 16'b0000010010110101;
            15'd15385: log10_cal = 16'b0000010010110101;
            15'd15386: log10_cal = 16'b0000010010110101;
            15'd15387: log10_cal = 16'b0000010010110101;
            15'd15388: log10_cal = 16'b0000010010110101;
            15'd15389: log10_cal = 16'b0000010010110101;
            15'd15390: log10_cal = 16'b0000010010110101;
            15'd15391: log10_cal = 16'b0000010010110101;
            15'd15392: log10_cal = 16'b0000010010110101;
            15'd15393: log10_cal = 16'b0000010010110101;
            15'd15394: log10_cal = 16'b0000010010110101;
            15'd15395: log10_cal = 16'b0000010010110101;
            15'd15396: log10_cal = 16'b0000010010110101;
            15'd15397: log10_cal = 16'b0000010010110101;
            15'd15398: log10_cal = 16'b0000010010110101;
            15'd15399: log10_cal = 16'b0000010010110101;
            15'd15400: log10_cal = 16'b0000010010110101;
            15'd15401: log10_cal = 16'b0000010010110101;
            15'd15402: log10_cal = 16'b0000010010110101;
            15'd15403: log10_cal = 16'b0000010010110101;
            15'd15404: log10_cal = 16'b0000010010110101;
            15'd15405: log10_cal = 16'b0000010010110101;
            15'd15406: log10_cal = 16'b0000010010110101;
            15'd15407: log10_cal = 16'b0000010010110101;
            15'd15408: log10_cal = 16'b0000010010110101;
            15'd15409: log10_cal = 16'b0000010010110101;
            15'd15410: log10_cal = 16'b0000010010110101;
            15'd15411: log10_cal = 16'b0000010010110101;
            15'd15412: log10_cal = 16'b0000010010110101;
            15'd15413: log10_cal = 16'b0000010010110101;
            15'd15414: log10_cal = 16'b0000010010110101;
            15'd15415: log10_cal = 16'b0000010010110101;
            15'd15416: log10_cal = 16'b0000010010110101;
            15'd15417: log10_cal = 16'b0000010010110101;
            15'd15418: log10_cal = 16'b0000010010110101;
            15'd15419: log10_cal = 16'b0000010010110110;
            15'd15420: log10_cal = 16'b0000010010110110;
            15'd15421: log10_cal = 16'b0000010010110110;
            15'd15422: log10_cal = 16'b0000010010110110;
            15'd15423: log10_cal = 16'b0000010010110110;
            15'd15424: log10_cal = 16'b0000010010110110;
            15'd15425: log10_cal = 16'b0000010010110110;
            15'd15426: log10_cal = 16'b0000010010110110;
            15'd15427: log10_cal = 16'b0000010010110110;
            15'd15428: log10_cal = 16'b0000010010110110;
            15'd15429: log10_cal = 16'b0000010010110110;
            15'd15430: log10_cal = 16'b0000010010110110;
            15'd15431: log10_cal = 16'b0000010010110110;
            15'd15432: log10_cal = 16'b0000010010110110;
            15'd15433: log10_cal = 16'b0000010010110110;
            15'd15434: log10_cal = 16'b0000010010110110;
            15'd15435: log10_cal = 16'b0000010010110110;
            15'd15436: log10_cal = 16'b0000010010110110;
            15'd15437: log10_cal = 16'b0000010010110110;
            15'd15438: log10_cal = 16'b0000010010110110;
            15'd15439: log10_cal = 16'b0000010010110110;
            15'd15440: log10_cal = 16'b0000010010110110;
            15'd15441: log10_cal = 16'b0000010010110110;
            15'd15442: log10_cal = 16'b0000010010110110;
            15'd15443: log10_cal = 16'b0000010010110110;
            15'd15444: log10_cal = 16'b0000010010110110;
            15'd15445: log10_cal = 16'b0000010010110110;
            15'd15446: log10_cal = 16'b0000010010110110;
            15'd15447: log10_cal = 16'b0000010010110110;
            15'd15448: log10_cal = 16'b0000010010110110;
            15'd15449: log10_cal = 16'b0000010010110110;
            15'd15450: log10_cal = 16'b0000010010110110;
            15'd15451: log10_cal = 16'b0000010010110110;
            15'd15452: log10_cal = 16'b0000010010110110;
            15'd15453: log10_cal = 16'b0000010010110111;
            15'd15454: log10_cal = 16'b0000010010110111;
            15'd15455: log10_cal = 16'b0000010010110111;
            15'd15456: log10_cal = 16'b0000010010110111;
            15'd15457: log10_cal = 16'b0000010010110111;
            15'd15458: log10_cal = 16'b0000010010110111;
            15'd15459: log10_cal = 16'b0000010010110111;
            15'd15460: log10_cal = 16'b0000010010110111;
            15'd15461: log10_cal = 16'b0000010010110111;
            15'd15462: log10_cal = 16'b0000010010110111;
            15'd15463: log10_cal = 16'b0000010010110111;
            15'd15464: log10_cal = 16'b0000010010110111;
            15'd15465: log10_cal = 16'b0000010010110111;
            15'd15466: log10_cal = 16'b0000010010110111;
            15'd15467: log10_cal = 16'b0000010010110111;
            15'd15468: log10_cal = 16'b0000010010110111;
            15'd15469: log10_cal = 16'b0000010010110111;
            15'd15470: log10_cal = 16'b0000010010110111;
            15'd15471: log10_cal = 16'b0000010010110111;
            15'd15472: log10_cal = 16'b0000010010110111;
            15'd15473: log10_cal = 16'b0000010010110111;
            15'd15474: log10_cal = 16'b0000010010110111;
            15'd15475: log10_cal = 16'b0000010010110111;
            15'd15476: log10_cal = 16'b0000010010110111;
            15'd15477: log10_cal = 16'b0000010010110111;
            15'd15478: log10_cal = 16'b0000010010110111;
            15'd15479: log10_cal = 16'b0000010010110111;
            15'd15480: log10_cal = 16'b0000010010110111;
            15'd15481: log10_cal = 16'b0000010010110111;
            15'd15482: log10_cal = 16'b0000010010110111;
            15'd15483: log10_cal = 16'b0000010010110111;
            15'd15484: log10_cal = 16'b0000010010110111;
            15'd15485: log10_cal = 16'b0000010010110111;
            15'd15486: log10_cal = 16'b0000010010110111;
            15'd15487: log10_cal = 16'b0000010010110111;
            15'd15488: log10_cal = 16'b0000010010111000;
            15'd15489: log10_cal = 16'b0000010010111000;
            15'd15490: log10_cal = 16'b0000010010111000;
            15'd15491: log10_cal = 16'b0000010010111000;
            15'd15492: log10_cal = 16'b0000010010111000;
            15'd15493: log10_cal = 16'b0000010010111000;
            15'd15494: log10_cal = 16'b0000010010111000;
            15'd15495: log10_cal = 16'b0000010010111000;
            15'd15496: log10_cal = 16'b0000010010111000;
            15'd15497: log10_cal = 16'b0000010010111000;
            15'd15498: log10_cal = 16'b0000010010111000;
            15'd15499: log10_cal = 16'b0000010010111000;
            15'd15500: log10_cal = 16'b0000010010111000;
            15'd15501: log10_cal = 16'b0000010010111000;
            15'd15502: log10_cal = 16'b0000010010111000;
            15'd15503: log10_cal = 16'b0000010010111000;
            15'd15504: log10_cal = 16'b0000010010111000;
            15'd15505: log10_cal = 16'b0000010010111000;
            15'd15506: log10_cal = 16'b0000010010111000;
            15'd15507: log10_cal = 16'b0000010010111000;
            15'd15508: log10_cal = 16'b0000010010111000;
            15'd15509: log10_cal = 16'b0000010010111000;
            15'd15510: log10_cal = 16'b0000010010111000;
            15'd15511: log10_cal = 16'b0000010010111000;
            15'd15512: log10_cal = 16'b0000010010111000;
            15'd15513: log10_cal = 16'b0000010010111000;
            15'd15514: log10_cal = 16'b0000010010111000;
            15'd15515: log10_cal = 16'b0000010010111000;
            15'd15516: log10_cal = 16'b0000010010111000;
            15'd15517: log10_cal = 16'b0000010010111000;
            15'd15518: log10_cal = 16'b0000010010111000;
            15'd15519: log10_cal = 16'b0000010010111000;
            15'd15520: log10_cal = 16'b0000010010111000;
            15'd15521: log10_cal = 16'b0000010010111000;
            15'd15522: log10_cal = 16'b0000010010111000;
            15'd15523: log10_cal = 16'b0000010010111001;
            15'd15524: log10_cal = 16'b0000010010111001;
            15'd15525: log10_cal = 16'b0000010010111001;
            15'd15526: log10_cal = 16'b0000010010111001;
            15'd15527: log10_cal = 16'b0000010010111001;
            15'd15528: log10_cal = 16'b0000010010111001;
            15'd15529: log10_cal = 16'b0000010010111001;
            15'd15530: log10_cal = 16'b0000010010111001;
            15'd15531: log10_cal = 16'b0000010010111001;
            15'd15532: log10_cal = 16'b0000010010111001;
            15'd15533: log10_cal = 16'b0000010010111001;
            15'd15534: log10_cal = 16'b0000010010111001;
            15'd15535: log10_cal = 16'b0000010010111001;
            15'd15536: log10_cal = 16'b0000010010111001;
            15'd15537: log10_cal = 16'b0000010010111001;
            15'd15538: log10_cal = 16'b0000010010111001;
            15'd15539: log10_cal = 16'b0000010010111001;
            15'd15540: log10_cal = 16'b0000010010111001;
            15'd15541: log10_cal = 16'b0000010010111001;
            15'd15542: log10_cal = 16'b0000010010111001;
            15'd15543: log10_cal = 16'b0000010010111001;
            15'd15544: log10_cal = 16'b0000010010111001;
            15'd15545: log10_cal = 16'b0000010010111001;
            15'd15546: log10_cal = 16'b0000010010111001;
            15'd15547: log10_cal = 16'b0000010010111001;
            15'd15548: log10_cal = 16'b0000010010111001;
            15'd15549: log10_cal = 16'b0000010010111001;
            15'd15550: log10_cal = 16'b0000010010111001;
            15'd15551: log10_cal = 16'b0000010010111001;
            15'd15552: log10_cal = 16'b0000010010111001;
            15'd15553: log10_cal = 16'b0000010010111001;
            15'd15554: log10_cal = 16'b0000010010111001;
            15'd15555: log10_cal = 16'b0000010010111001;
            15'd15556: log10_cal = 16'b0000010010111001;
            15'd15557: log10_cal = 16'b0000010010111001;
            15'd15558: log10_cal = 16'b0000010010111010;
            15'd15559: log10_cal = 16'b0000010010111010;
            15'd15560: log10_cal = 16'b0000010010111010;
            15'd15561: log10_cal = 16'b0000010010111010;
            15'd15562: log10_cal = 16'b0000010010111010;
            15'd15563: log10_cal = 16'b0000010010111010;
            15'd15564: log10_cal = 16'b0000010010111010;
            15'd15565: log10_cal = 16'b0000010010111010;
            15'd15566: log10_cal = 16'b0000010010111010;
            15'd15567: log10_cal = 16'b0000010010111010;
            15'd15568: log10_cal = 16'b0000010010111010;
            15'd15569: log10_cal = 16'b0000010010111010;
            15'd15570: log10_cal = 16'b0000010010111010;
            15'd15571: log10_cal = 16'b0000010010111010;
            15'd15572: log10_cal = 16'b0000010010111010;
            15'd15573: log10_cal = 16'b0000010010111010;
            15'd15574: log10_cal = 16'b0000010010111010;
            15'd15575: log10_cal = 16'b0000010010111010;
            15'd15576: log10_cal = 16'b0000010010111010;
            15'd15577: log10_cal = 16'b0000010010111010;
            15'd15578: log10_cal = 16'b0000010010111010;
            15'd15579: log10_cal = 16'b0000010010111010;
            15'd15580: log10_cal = 16'b0000010010111010;
            15'd15581: log10_cal = 16'b0000010010111010;
            15'd15582: log10_cal = 16'b0000010010111010;
            15'd15583: log10_cal = 16'b0000010010111010;
            15'd15584: log10_cal = 16'b0000010010111010;
            15'd15585: log10_cal = 16'b0000010010111010;
            15'd15586: log10_cal = 16'b0000010010111010;
            15'd15587: log10_cal = 16'b0000010010111010;
            15'd15588: log10_cal = 16'b0000010010111010;
            15'd15589: log10_cal = 16'b0000010010111010;
            15'd15590: log10_cal = 16'b0000010010111010;
            15'd15591: log10_cal = 16'b0000010010111010;
            15'd15592: log10_cal = 16'b0000010010111010;
            15'd15593: log10_cal = 16'b0000010010111011;
            15'd15594: log10_cal = 16'b0000010010111011;
            15'd15595: log10_cal = 16'b0000010010111011;
            15'd15596: log10_cal = 16'b0000010010111011;
            15'd15597: log10_cal = 16'b0000010010111011;
            15'd15598: log10_cal = 16'b0000010010111011;
            15'd15599: log10_cal = 16'b0000010010111011;
            15'd15600: log10_cal = 16'b0000010010111011;
            15'd15601: log10_cal = 16'b0000010010111011;
            15'd15602: log10_cal = 16'b0000010010111011;
            15'd15603: log10_cal = 16'b0000010010111011;
            15'd15604: log10_cal = 16'b0000010010111011;
            15'd15605: log10_cal = 16'b0000010010111011;
            15'd15606: log10_cal = 16'b0000010010111011;
            15'd15607: log10_cal = 16'b0000010010111011;
            15'd15608: log10_cal = 16'b0000010010111011;
            15'd15609: log10_cal = 16'b0000010010111011;
            15'd15610: log10_cal = 16'b0000010010111011;
            15'd15611: log10_cal = 16'b0000010010111011;
            15'd15612: log10_cal = 16'b0000010010111011;
            15'd15613: log10_cal = 16'b0000010010111011;
            15'd15614: log10_cal = 16'b0000010010111011;
            15'd15615: log10_cal = 16'b0000010010111011;
            15'd15616: log10_cal = 16'b0000010010111011;
            15'd15617: log10_cal = 16'b0000010010111011;
            15'd15618: log10_cal = 16'b0000010010111011;
            15'd15619: log10_cal = 16'b0000010010111011;
            15'd15620: log10_cal = 16'b0000010010111011;
            15'd15621: log10_cal = 16'b0000010010111011;
            15'd15622: log10_cal = 16'b0000010010111011;
            15'd15623: log10_cal = 16'b0000010010111011;
            15'd15624: log10_cal = 16'b0000010010111011;
            15'd15625: log10_cal = 16'b0000010010111011;
            15'd15626: log10_cal = 16'b0000010010111011;
            15'd15627: log10_cal = 16'b0000010010111011;
            15'd15628: log10_cal = 16'b0000010010111100;
            15'd15629: log10_cal = 16'b0000010010111100;
            15'd15630: log10_cal = 16'b0000010010111100;
            15'd15631: log10_cal = 16'b0000010010111100;
            15'd15632: log10_cal = 16'b0000010010111100;
            15'd15633: log10_cal = 16'b0000010010111100;
            15'd15634: log10_cal = 16'b0000010010111100;
            15'd15635: log10_cal = 16'b0000010010111100;
            15'd15636: log10_cal = 16'b0000010010111100;
            15'd15637: log10_cal = 16'b0000010010111100;
            15'd15638: log10_cal = 16'b0000010010111100;
            15'd15639: log10_cal = 16'b0000010010111100;
            15'd15640: log10_cal = 16'b0000010010111100;
            15'd15641: log10_cal = 16'b0000010010111100;
            15'd15642: log10_cal = 16'b0000010010111100;
            15'd15643: log10_cal = 16'b0000010010111100;
            15'd15644: log10_cal = 16'b0000010010111100;
            15'd15645: log10_cal = 16'b0000010010111100;
            15'd15646: log10_cal = 16'b0000010010111100;
            15'd15647: log10_cal = 16'b0000010010111100;
            15'd15648: log10_cal = 16'b0000010010111100;
            15'd15649: log10_cal = 16'b0000010010111100;
            15'd15650: log10_cal = 16'b0000010010111100;
            15'd15651: log10_cal = 16'b0000010010111100;
            15'd15652: log10_cal = 16'b0000010010111100;
            15'd15653: log10_cal = 16'b0000010010111100;
            15'd15654: log10_cal = 16'b0000010010111100;
            15'd15655: log10_cal = 16'b0000010010111100;
            15'd15656: log10_cal = 16'b0000010010111100;
            15'd15657: log10_cal = 16'b0000010010111100;
            15'd15658: log10_cal = 16'b0000010010111100;
            15'd15659: log10_cal = 16'b0000010010111100;
            15'd15660: log10_cal = 16'b0000010010111100;
            15'd15661: log10_cal = 16'b0000010010111100;
            15'd15662: log10_cal = 16'b0000010010111100;
            15'd15663: log10_cal = 16'b0000010010111101;
            15'd15664: log10_cal = 16'b0000010010111101;
            15'd15665: log10_cal = 16'b0000010010111101;
            15'd15666: log10_cal = 16'b0000010010111101;
            15'd15667: log10_cal = 16'b0000010010111101;
            15'd15668: log10_cal = 16'b0000010010111101;
            15'd15669: log10_cal = 16'b0000010010111101;
            15'd15670: log10_cal = 16'b0000010010111101;
            15'd15671: log10_cal = 16'b0000010010111101;
            15'd15672: log10_cal = 16'b0000010010111101;
            15'd15673: log10_cal = 16'b0000010010111101;
            15'd15674: log10_cal = 16'b0000010010111101;
            15'd15675: log10_cal = 16'b0000010010111101;
            15'd15676: log10_cal = 16'b0000010010111101;
            15'd15677: log10_cal = 16'b0000010010111101;
            15'd15678: log10_cal = 16'b0000010010111101;
            15'd15679: log10_cal = 16'b0000010010111101;
            15'd15680: log10_cal = 16'b0000010010111101;
            15'd15681: log10_cal = 16'b0000010010111101;
            15'd15682: log10_cal = 16'b0000010010111101;
            15'd15683: log10_cal = 16'b0000010010111101;
            15'd15684: log10_cal = 16'b0000010010111101;
            15'd15685: log10_cal = 16'b0000010010111101;
            15'd15686: log10_cal = 16'b0000010010111101;
            15'd15687: log10_cal = 16'b0000010010111101;
            15'd15688: log10_cal = 16'b0000010010111101;
            15'd15689: log10_cal = 16'b0000010010111101;
            15'd15690: log10_cal = 16'b0000010010111101;
            15'd15691: log10_cal = 16'b0000010010111101;
            15'd15692: log10_cal = 16'b0000010010111101;
            15'd15693: log10_cal = 16'b0000010010111101;
            15'd15694: log10_cal = 16'b0000010010111101;
            15'd15695: log10_cal = 16'b0000010010111101;
            15'd15696: log10_cal = 16'b0000010010111101;
            15'd15697: log10_cal = 16'b0000010010111101;
            15'd15698: log10_cal = 16'b0000010010111101;
            15'd15699: log10_cal = 16'b0000010010111110;
            15'd15700: log10_cal = 16'b0000010010111110;
            15'd15701: log10_cal = 16'b0000010010111110;
            15'd15702: log10_cal = 16'b0000010010111110;
            15'd15703: log10_cal = 16'b0000010010111110;
            15'd15704: log10_cal = 16'b0000010010111110;
            15'd15705: log10_cal = 16'b0000010010111110;
            15'd15706: log10_cal = 16'b0000010010111110;
            15'd15707: log10_cal = 16'b0000010010111110;
            15'd15708: log10_cal = 16'b0000010010111110;
            15'd15709: log10_cal = 16'b0000010010111110;
            15'd15710: log10_cal = 16'b0000010010111110;
            15'd15711: log10_cal = 16'b0000010010111110;
            15'd15712: log10_cal = 16'b0000010010111110;
            15'd15713: log10_cal = 16'b0000010010111110;
            15'd15714: log10_cal = 16'b0000010010111110;
            15'd15715: log10_cal = 16'b0000010010111110;
            15'd15716: log10_cal = 16'b0000010010111110;
            15'd15717: log10_cal = 16'b0000010010111110;
            15'd15718: log10_cal = 16'b0000010010111110;
            15'd15719: log10_cal = 16'b0000010010111110;
            15'd15720: log10_cal = 16'b0000010010111110;
            15'd15721: log10_cal = 16'b0000010010111110;
            15'd15722: log10_cal = 16'b0000010010111110;
            15'd15723: log10_cal = 16'b0000010010111110;
            15'd15724: log10_cal = 16'b0000010010111110;
            15'd15725: log10_cal = 16'b0000010010111110;
            15'd15726: log10_cal = 16'b0000010010111110;
            15'd15727: log10_cal = 16'b0000010010111110;
            15'd15728: log10_cal = 16'b0000010010111110;
            15'd15729: log10_cal = 16'b0000010010111110;
            15'd15730: log10_cal = 16'b0000010010111110;
            15'd15731: log10_cal = 16'b0000010010111110;
            15'd15732: log10_cal = 16'b0000010010111110;
            15'd15733: log10_cal = 16'b0000010010111110;
            15'd15734: log10_cal = 16'b0000010010111111;
            15'd15735: log10_cal = 16'b0000010010111111;
            15'd15736: log10_cal = 16'b0000010010111111;
            15'd15737: log10_cal = 16'b0000010010111111;
            15'd15738: log10_cal = 16'b0000010010111111;
            15'd15739: log10_cal = 16'b0000010010111111;
            15'd15740: log10_cal = 16'b0000010010111111;
            15'd15741: log10_cal = 16'b0000010010111111;
            15'd15742: log10_cal = 16'b0000010010111111;
            15'd15743: log10_cal = 16'b0000010010111111;
            15'd15744: log10_cal = 16'b0000010010111111;
            15'd15745: log10_cal = 16'b0000010010111111;
            15'd15746: log10_cal = 16'b0000010010111111;
            15'd15747: log10_cal = 16'b0000010010111111;
            15'd15748: log10_cal = 16'b0000010010111111;
            15'd15749: log10_cal = 16'b0000010010111111;
            15'd15750: log10_cal = 16'b0000010010111111;
            15'd15751: log10_cal = 16'b0000010010111111;
            15'd15752: log10_cal = 16'b0000010010111111;
            15'd15753: log10_cal = 16'b0000010010111111;
            15'd15754: log10_cal = 16'b0000010010111111;
            15'd15755: log10_cal = 16'b0000010010111111;
            15'd15756: log10_cal = 16'b0000010010111111;
            15'd15757: log10_cal = 16'b0000010010111111;
            15'd15758: log10_cal = 16'b0000010010111111;
            15'd15759: log10_cal = 16'b0000010010111111;
            15'd15760: log10_cal = 16'b0000010010111111;
            15'd15761: log10_cal = 16'b0000010010111111;
            15'd15762: log10_cal = 16'b0000010010111111;
            15'd15763: log10_cal = 16'b0000010010111111;
            15'd15764: log10_cal = 16'b0000010010111111;
            15'd15765: log10_cal = 16'b0000010010111111;
            15'd15766: log10_cal = 16'b0000010010111111;
            15'd15767: log10_cal = 16'b0000010010111111;
            15'd15768: log10_cal = 16'b0000010010111111;
            15'd15769: log10_cal = 16'b0000010011000000;
            15'd15770: log10_cal = 16'b0000010011000000;
            15'd15771: log10_cal = 16'b0000010011000000;
            15'd15772: log10_cal = 16'b0000010011000000;
            15'd15773: log10_cal = 16'b0000010011000000;
            15'd15774: log10_cal = 16'b0000010011000000;
            15'd15775: log10_cal = 16'b0000010011000000;
            15'd15776: log10_cal = 16'b0000010011000000;
            15'd15777: log10_cal = 16'b0000010011000000;
            15'd15778: log10_cal = 16'b0000010011000000;
            15'd15779: log10_cal = 16'b0000010011000000;
            15'd15780: log10_cal = 16'b0000010011000000;
            15'd15781: log10_cal = 16'b0000010011000000;
            15'd15782: log10_cal = 16'b0000010011000000;
            15'd15783: log10_cal = 16'b0000010011000000;
            15'd15784: log10_cal = 16'b0000010011000000;
            15'd15785: log10_cal = 16'b0000010011000000;
            15'd15786: log10_cal = 16'b0000010011000000;
            15'd15787: log10_cal = 16'b0000010011000000;
            15'd15788: log10_cal = 16'b0000010011000000;
            15'd15789: log10_cal = 16'b0000010011000000;
            15'd15790: log10_cal = 16'b0000010011000000;
            15'd15791: log10_cal = 16'b0000010011000000;
            15'd15792: log10_cal = 16'b0000010011000000;
            15'd15793: log10_cal = 16'b0000010011000000;
            15'd15794: log10_cal = 16'b0000010011000000;
            15'd15795: log10_cal = 16'b0000010011000000;
            15'd15796: log10_cal = 16'b0000010011000000;
            15'd15797: log10_cal = 16'b0000010011000000;
            15'd15798: log10_cal = 16'b0000010011000000;
            15'd15799: log10_cal = 16'b0000010011000000;
            15'd15800: log10_cal = 16'b0000010011000000;
            15'd15801: log10_cal = 16'b0000010011000000;
            15'd15802: log10_cal = 16'b0000010011000000;
            15'd15803: log10_cal = 16'b0000010011000000;
            15'd15804: log10_cal = 16'b0000010011000000;
            15'd15805: log10_cal = 16'b0000010011000001;
            15'd15806: log10_cal = 16'b0000010011000001;
            15'd15807: log10_cal = 16'b0000010011000001;
            15'd15808: log10_cal = 16'b0000010011000001;
            15'd15809: log10_cal = 16'b0000010011000001;
            15'd15810: log10_cal = 16'b0000010011000001;
            15'd15811: log10_cal = 16'b0000010011000001;
            15'd15812: log10_cal = 16'b0000010011000001;
            15'd15813: log10_cal = 16'b0000010011000001;
            15'd15814: log10_cal = 16'b0000010011000001;
            15'd15815: log10_cal = 16'b0000010011000001;
            15'd15816: log10_cal = 16'b0000010011000001;
            15'd15817: log10_cal = 16'b0000010011000001;
            15'd15818: log10_cal = 16'b0000010011000001;
            15'd15819: log10_cal = 16'b0000010011000001;
            15'd15820: log10_cal = 16'b0000010011000001;
            15'd15821: log10_cal = 16'b0000010011000001;
            15'd15822: log10_cal = 16'b0000010011000001;
            15'd15823: log10_cal = 16'b0000010011000001;
            15'd15824: log10_cal = 16'b0000010011000001;
            15'd15825: log10_cal = 16'b0000010011000001;
            15'd15826: log10_cal = 16'b0000010011000001;
            15'd15827: log10_cal = 16'b0000010011000001;
            15'd15828: log10_cal = 16'b0000010011000001;
            15'd15829: log10_cal = 16'b0000010011000001;
            15'd15830: log10_cal = 16'b0000010011000001;
            15'd15831: log10_cal = 16'b0000010011000001;
            15'd15832: log10_cal = 16'b0000010011000001;
            15'd15833: log10_cal = 16'b0000010011000001;
            15'd15834: log10_cal = 16'b0000010011000001;
            15'd15835: log10_cal = 16'b0000010011000001;
            15'd15836: log10_cal = 16'b0000010011000001;
            15'd15837: log10_cal = 16'b0000010011000001;
            15'd15838: log10_cal = 16'b0000010011000001;
            15'd15839: log10_cal = 16'b0000010011000001;
            15'd15840: log10_cal = 16'b0000010011000010;
            15'd15841: log10_cal = 16'b0000010011000010;
            15'd15842: log10_cal = 16'b0000010011000010;
            15'd15843: log10_cal = 16'b0000010011000010;
            15'd15844: log10_cal = 16'b0000010011000010;
            15'd15845: log10_cal = 16'b0000010011000010;
            15'd15846: log10_cal = 16'b0000010011000010;
            15'd15847: log10_cal = 16'b0000010011000010;
            15'd15848: log10_cal = 16'b0000010011000010;
            15'd15849: log10_cal = 16'b0000010011000010;
            15'd15850: log10_cal = 16'b0000010011000010;
            15'd15851: log10_cal = 16'b0000010011000010;
            15'd15852: log10_cal = 16'b0000010011000010;
            15'd15853: log10_cal = 16'b0000010011000010;
            15'd15854: log10_cal = 16'b0000010011000010;
            15'd15855: log10_cal = 16'b0000010011000010;
            15'd15856: log10_cal = 16'b0000010011000010;
            15'd15857: log10_cal = 16'b0000010011000010;
            15'd15858: log10_cal = 16'b0000010011000010;
            15'd15859: log10_cal = 16'b0000010011000010;
            15'd15860: log10_cal = 16'b0000010011000010;
            15'd15861: log10_cal = 16'b0000010011000010;
            15'd15862: log10_cal = 16'b0000010011000010;
            15'd15863: log10_cal = 16'b0000010011000010;
            15'd15864: log10_cal = 16'b0000010011000010;
            15'd15865: log10_cal = 16'b0000010011000010;
            15'd15866: log10_cal = 16'b0000010011000010;
            15'd15867: log10_cal = 16'b0000010011000010;
            15'd15868: log10_cal = 16'b0000010011000010;
            15'd15869: log10_cal = 16'b0000010011000010;
            15'd15870: log10_cal = 16'b0000010011000010;
            15'd15871: log10_cal = 16'b0000010011000010;
            15'd15872: log10_cal = 16'b0000010011000010;
            15'd15873: log10_cal = 16'b0000010011000010;
            15'd15874: log10_cal = 16'b0000010011000010;
            15'd15875: log10_cal = 16'b0000010011000010;
            15'd15876: log10_cal = 16'b0000010011000011;
            15'd15877: log10_cal = 16'b0000010011000011;
            15'd15878: log10_cal = 16'b0000010011000011;
            15'd15879: log10_cal = 16'b0000010011000011;
            15'd15880: log10_cal = 16'b0000010011000011;
            15'd15881: log10_cal = 16'b0000010011000011;
            15'd15882: log10_cal = 16'b0000010011000011;
            15'd15883: log10_cal = 16'b0000010011000011;
            15'd15884: log10_cal = 16'b0000010011000011;
            15'd15885: log10_cal = 16'b0000010011000011;
            15'd15886: log10_cal = 16'b0000010011000011;
            15'd15887: log10_cal = 16'b0000010011000011;
            15'd15888: log10_cal = 16'b0000010011000011;
            15'd15889: log10_cal = 16'b0000010011000011;
            15'd15890: log10_cal = 16'b0000010011000011;
            15'd15891: log10_cal = 16'b0000010011000011;
            15'd15892: log10_cal = 16'b0000010011000011;
            15'd15893: log10_cal = 16'b0000010011000011;
            15'd15894: log10_cal = 16'b0000010011000011;
            15'd15895: log10_cal = 16'b0000010011000011;
            15'd15896: log10_cal = 16'b0000010011000011;
            15'd15897: log10_cal = 16'b0000010011000011;
            15'd15898: log10_cal = 16'b0000010011000011;
            15'd15899: log10_cal = 16'b0000010011000011;
            15'd15900: log10_cal = 16'b0000010011000011;
            15'd15901: log10_cal = 16'b0000010011000011;
            15'd15902: log10_cal = 16'b0000010011000011;
            15'd15903: log10_cal = 16'b0000010011000011;
            15'd15904: log10_cal = 16'b0000010011000011;
            15'd15905: log10_cal = 16'b0000010011000011;
            15'd15906: log10_cal = 16'b0000010011000011;
            15'd15907: log10_cal = 16'b0000010011000011;
            15'd15908: log10_cal = 16'b0000010011000011;
            15'd15909: log10_cal = 16'b0000010011000011;
            15'd15910: log10_cal = 16'b0000010011000011;
            15'd15911: log10_cal = 16'b0000010011000011;
            15'd15912: log10_cal = 16'b0000010011000100;
            15'd15913: log10_cal = 16'b0000010011000100;
            15'd15914: log10_cal = 16'b0000010011000100;
            15'd15915: log10_cal = 16'b0000010011000100;
            15'd15916: log10_cal = 16'b0000010011000100;
            15'd15917: log10_cal = 16'b0000010011000100;
            15'd15918: log10_cal = 16'b0000010011000100;
            15'd15919: log10_cal = 16'b0000010011000100;
            15'd15920: log10_cal = 16'b0000010011000100;
            15'd15921: log10_cal = 16'b0000010011000100;
            15'd15922: log10_cal = 16'b0000010011000100;
            15'd15923: log10_cal = 16'b0000010011000100;
            15'd15924: log10_cal = 16'b0000010011000100;
            15'd15925: log10_cal = 16'b0000010011000100;
            15'd15926: log10_cal = 16'b0000010011000100;
            15'd15927: log10_cal = 16'b0000010011000100;
            15'd15928: log10_cal = 16'b0000010011000100;
            15'd15929: log10_cal = 16'b0000010011000100;
            15'd15930: log10_cal = 16'b0000010011000100;
            15'd15931: log10_cal = 16'b0000010011000100;
            15'd15932: log10_cal = 16'b0000010011000100;
            15'd15933: log10_cal = 16'b0000010011000100;
            15'd15934: log10_cal = 16'b0000010011000100;
            15'd15935: log10_cal = 16'b0000010011000100;
            15'd15936: log10_cal = 16'b0000010011000100;
            15'd15937: log10_cal = 16'b0000010011000100;
            15'd15938: log10_cal = 16'b0000010011000100;
            15'd15939: log10_cal = 16'b0000010011000100;
            15'd15940: log10_cal = 16'b0000010011000100;
            15'd15941: log10_cal = 16'b0000010011000100;
            15'd15942: log10_cal = 16'b0000010011000100;
            15'd15943: log10_cal = 16'b0000010011000100;
            15'd15944: log10_cal = 16'b0000010011000100;
            15'd15945: log10_cal = 16'b0000010011000100;
            15'd15946: log10_cal = 16'b0000010011000100;
            15'd15947: log10_cal = 16'b0000010011000100;
            15'd15948: log10_cal = 16'b0000010011000101;
            15'd15949: log10_cal = 16'b0000010011000101;
            15'd15950: log10_cal = 16'b0000010011000101;
            15'd15951: log10_cal = 16'b0000010011000101;
            15'd15952: log10_cal = 16'b0000010011000101;
            15'd15953: log10_cal = 16'b0000010011000101;
            15'd15954: log10_cal = 16'b0000010011000101;
            15'd15955: log10_cal = 16'b0000010011000101;
            15'd15956: log10_cal = 16'b0000010011000101;
            15'd15957: log10_cal = 16'b0000010011000101;
            15'd15958: log10_cal = 16'b0000010011000101;
            15'd15959: log10_cal = 16'b0000010011000101;
            15'd15960: log10_cal = 16'b0000010011000101;
            15'd15961: log10_cal = 16'b0000010011000101;
            15'd15962: log10_cal = 16'b0000010011000101;
            15'd15963: log10_cal = 16'b0000010011000101;
            15'd15964: log10_cal = 16'b0000010011000101;
            15'd15965: log10_cal = 16'b0000010011000101;
            15'd15966: log10_cal = 16'b0000010011000101;
            15'd15967: log10_cal = 16'b0000010011000101;
            15'd15968: log10_cal = 16'b0000010011000101;
            15'd15969: log10_cal = 16'b0000010011000101;
            15'd15970: log10_cal = 16'b0000010011000101;
            15'd15971: log10_cal = 16'b0000010011000101;
            15'd15972: log10_cal = 16'b0000010011000101;
            15'd15973: log10_cal = 16'b0000010011000101;
            15'd15974: log10_cal = 16'b0000010011000101;
            15'd15975: log10_cal = 16'b0000010011000101;
            15'd15976: log10_cal = 16'b0000010011000101;
            15'd15977: log10_cal = 16'b0000010011000101;
            15'd15978: log10_cal = 16'b0000010011000101;
            15'd15979: log10_cal = 16'b0000010011000101;
            15'd15980: log10_cal = 16'b0000010011000101;
            15'd15981: log10_cal = 16'b0000010011000101;
            15'd15982: log10_cal = 16'b0000010011000101;
            15'd15983: log10_cal = 16'b0000010011000101;
            15'd15984: log10_cal = 16'b0000010011000110;
            15'd15985: log10_cal = 16'b0000010011000110;
            15'd15986: log10_cal = 16'b0000010011000110;
            15'd15987: log10_cal = 16'b0000010011000110;
            15'd15988: log10_cal = 16'b0000010011000110;
            15'd15989: log10_cal = 16'b0000010011000110;
            15'd15990: log10_cal = 16'b0000010011000110;
            15'd15991: log10_cal = 16'b0000010011000110;
            15'd15992: log10_cal = 16'b0000010011000110;
            15'd15993: log10_cal = 16'b0000010011000110;
            15'd15994: log10_cal = 16'b0000010011000110;
            15'd15995: log10_cal = 16'b0000010011000110;
            15'd15996: log10_cal = 16'b0000010011000110;
            15'd15997: log10_cal = 16'b0000010011000110;
            15'd15998: log10_cal = 16'b0000010011000110;
            15'd15999: log10_cal = 16'b0000010011000110;
            15'd16000: log10_cal = 16'b0000010011000110;
            15'd16001: log10_cal = 16'b0000010011000110;
            15'd16002: log10_cal = 16'b0000010011000110;
            15'd16003: log10_cal = 16'b0000010011000110;
            15'd16004: log10_cal = 16'b0000010011000110;
            15'd16005: log10_cal = 16'b0000010011000110;
            15'd16006: log10_cal = 16'b0000010011000110;
            15'd16007: log10_cal = 16'b0000010011000110;
            15'd16008: log10_cal = 16'b0000010011000110;
            15'd16009: log10_cal = 16'b0000010011000110;
            15'd16010: log10_cal = 16'b0000010011000110;
            15'd16011: log10_cal = 16'b0000010011000110;
            15'd16012: log10_cal = 16'b0000010011000110;
            15'd16013: log10_cal = 16'b0000010011000110;
            15'd16014: log10_cal = 16'b0000010011000110;
            15'd16015: log10_cal = 16'b0000010011000110;
            15'd16016: log10_cal = 16'b0000010011000110;
            15'd16017: log10_cal = 16'b0000010011000110;
            15'd16018: log10_cal = 16'b0000010011000110;
            15'd16019: log10_cal = 16'b0000010011000110;
            15'd16020: log10_cal = 16'b0000010011000111;
            15'd16021: log10_cal = 16'b0000010011000111;
            15'd16022: log10_cal = 16'b0000010011000111;
            15'd16023: log10_cal = 16'b0000010011000111;
            15'd16024: log10_cal = 16'b0000010011000111;
            15'd16025: log10_cal = 16'b0000010011000111;
            15'd16026: log10_cal = 16'b0000010011000111;
            15'd16027: log10_cal = 16'b0000010011000111;
            15'd16028: log10_cal = 16'b0000010011000111;
            15'd16029: log10_cal = 16'b0000010011000111;
            15'd16030: log10_cal = 16'b0000010011000111;
            15'd16031: log10_cal = 16'b0000010011000111;
            15'd16032: log10_cal = 16'b0000010011000111;
            15'd16033: log10_cal = 16'b0000010011000111;
            15'd16034: log10_cal = 16'b0000010011000111;
            15'd16035: log10_cal = 16'b0000010011000111;
            15'd16036: log10_cal = 16'b0000010011000111;
            15'd16037: log10_cal = 16'b0000010011000111;
            15'd16038: log10_cal = 16'b0000010011000111;
            15'd16039: log10_cal = 16'b0000010011000111;
            15'd16040: log10_cal = 16'b0000010011000111;
            15'd16041: log10_cal = 16'b0000010011000111;
            15'd16042: log10_cal = 16'b0000010011000111;
            15'd16043: log10_cal = 16'b0000010011000111;
            15'd16044: log10_cal = 16'b0000010011000111;
            15'd16045: log10_cal = 16'b0000010011000111;
            15'd16046: log10_cal = 16'b0000010011000111;
            15'd16047: log10_cal = 16'b0000010011000111;
            15'd16048: log10_cal = 16'b0000010011000111;
            15'd16049: log10_cal = 16'b0000010011000111;
            15'd16050: log10_cal = 16'b0000010011000111;
            15'd16051: log10_cal = 16'b0000010011000111;
            15'd16052: log10_cal = 16'b0000010011000111;
            15'd16053: log10_cal = 16'b0000010011000111;
            15'd16054: log10_cal = 16'b0000010011000111;
            15'd16055: log10_cal = 16'b0000010011000111;
            15'd16056: log10_cal = 16'b0000010011001000;
            15'd16057: log10_cal = 16'b0000010011001000;
            15'd16058: log10_cal = 16'b0000010011001000;
            15'd16059: log10_cal = 16'b0000010011001000;
            15'd16060: log10_cal = 16'b0000010011001000;
            15'd16061: log10_cal = 16'b0000010011001000;
            15'd16062: log10_cal = 16'b0000010011001000;
            15'd16063: log10_cal = 16'b0000010011001000;
            15'd16064: log10_cal = 16'b0000010011001000;
            15'd16065: log10_cal = 16'b0000010011001000;
            15'd16066: log10_cal = 16'b0000010011001000;
            15'd16067: log10_cal = 16'b0000010011001000;
            15'd16068: log10_cal = 16'b0000010011001000;
            15'd16069: log10_cal = 16'b0000010011001000;
            15'd16070: log10_cal = 16'b0000010011001000;
            15'd16071: log10_cal = 16'b0000010011001000;
            15'd16072: log10_cal = 16'b0000010011001000;
            15'd16073: log10_cal = 16'b0000010011001000;
            15'd16074: log10_cal = 16'b0000010011001000;
            15'd16075: log10_cal = 16'b0000010011001000;
            15'd16076: log10_cal = 16'b0000010011001000;
            15'd16077: log10_cal = 16'b0000010011001000;
            15'd16078: log10_cal = 16'b0000010011001000;
            15'd16079: log10_cal = 16'b0000010011001000;
            15'd16080: log10_cal = 16'b0000010011001000;
            15'd16081: log10_cal = 16'b0000010011001000;
            15'd16082: log10_cal = 16'b0000010011001000;
            15'd16083: log10_cal = 16'b0000010011001000;
            15'd16084: log10_cal = 16'b0000010011001000;
            15'd16085: log10_cal = 16'b0000010011001000;
            15'd16086: log10_cal = 16'b0000010011001000;
            15'd16087: log10_cal = 16'b0000010011001000;
            15'd16088: log10_cal = 16'b0000010011001000;
            15'd16089: log10_cal = 16'b0000010011001000;
            15'd16090: log10_cal = 16'b0000010011001000;
            15'd16091: log10_cal = 16'b0000010011001000;
            15'd16092: log10_cal = 16'b0000010011001001;
            15'd16093: log10_cal = 16'b0000010011001001;
            15'd16094: log10_cal = 16'b0000010011001001;
            15'd16095: log10_cal = 16'b0000010011001001;
            15'd16096: log10_cal = 16'b0000010011001001;
            15'd16097: log10_cal = 16'b0000010011001001;
            15'd16098: log10_cal = 16'b0000010011001001;
            15'd16099: log10_cal = 16'b0000010011001001;
            15'd16100: log10_cal = 16'b0000010011001001;
            15'd16101: log10_cal = 16'b0000010011001001;
            15'd16102: log10_cal = 16'b0000010011001001;
            15'd16103: log10_cal = 16'b0000010011001001;
            15'd16104: log10_cal = 16'b0000010011001001;
            15'd16105: log10_cal = 16'b0000010011001001;
            15'd16106: log10_cal = 16'b0000010011001001;
            15'd16107: log10_cal = 16'b0000010011001001;
            15'd16108: log10_cal = 16'b0000010011001001;
            15'd16109: log10_cal = 16'b0000010011001001;
            15'd16110: log10_cal = 16'b0000010011001001;
            15'd16111: log10_cal = 16'b0000010011001001;
            15'd16112: log10_cal = 16'b0000010011001001;
            15'd16113: log10_cal = 16'b0000010011001001;
            15'd16114: log10_cal = 16'b0000010011001001;
            15'd16115: log10_cal = 16'b0000010011001001;
            15'd16116: log10_cal = 16'b0000010011001001;
            15'd16117: log10_cal = 16'b0000010011001001;
            15'd16118: log10_cal = 16'b0000010011001001;
            15'd16119: log10_cal = 16'b0000010011001001;
            15'd16120: log10_cal = 16'b0000010011001001;
            15'd16121: log10_cal = 16'b0000010011001001;
            15'd16122: log10_cal = 16'b0000010011001001;
            15'd16123: log10_cal = 16'b0000010011001001;
            15'd16124: log10_cal = 16'b0000010011001001;
            15'd16125: log10_cal = 16'b0000010011001001;
            15'd16126: log10_cal = 16'b0000010011001001;
            15'd16127: log10_cal = 16'b0000010011001001;
            15'd16128: log10_cal = 16'b0000010011001010;
            15'd16129: log10_cal = 16'b0000010011001010;
            15'd16130: log10_cal = 16'b0000010011001010;
            15'd16131: log10_cal = 16'b0000010011001010;
            15'd16132: log10_cal = 16'b0000010011001010;
            15'd16133: log10_cal = 16'b0000010011001010;
            15'd16134: log10_cal = 16'b0000010011001010;
            15'd16135: log10_cal = 16'b0000010011001010;
            15'd16136: log10_cal = 16'b0000010011001010;
            15'd16137: log10_cal = 16'b0000010011001010;
            15'd16138: log10_cal = 16'b0000010011001010;
            15'd16139: log10_cal = 16'b0000010011001010;
            15'd16140: log10_cal = 16'b0000010011001010;
            15'd16141: log10_cal = 16'b0000010011001010;
            15'd16142: log10_cal = 16'b0000010011001010;
            15'd16143: log10_cal = 16'b0000010011001010;
            15'd16144: log10_cal = 16'b0000010011001010;
            15'd16145: log10_cal = 16'b0000010011001010;
            15'd16146: log10_cal = 16'b0000010011001010;
            15'd16147: log10_cal = 16'b0000010011001010;
            15'd16148: log10_cal = 16'b0000010011001010;
            15'd16149: log10_cal = 16'b0000010011001010;
            15'd16150: log10_cal = 16'b0000010011001010;
            15'd16151: log10_cal = 16'b0000010011001010;
            15'd16152: log10_cal = 16'b0000010011001010;
            15'd16153: log10_cal = 16'b0000010011001010;
            15'd16154: log10_cal = 16'b0000010011001010;
            15'd16155: log10_cal = 16'b0000010011001010;
            15'd16156: log10_cal = 16'b0000010011001010;
            15'd16157: log10_cal = 16'b0000010011001010;
            15'd16158: log10_cal = 16'b0000010011001010;
            15'd16159: log10_cal = 16'b0000010011001010;
            15'd16160: log10_cal = 16'b0000010011001010;
            15'd16161: log10_cal = 16'b0000010011001010;
            15'd16162: log10_cal = 16'b0000010011001010;
            15'd16163: log10_cal = 16'b0000010011001010;
            15'd16164: log10_cal = 16'b0000010011001011;
            15'd16165: log10_cal = 16'b0000010011001011;
            15'd16166: log10_cal = 16'b0000010011001011;
            15'd16167: log10_cal = 16'b0000010011001011;
            15'd16168: log10_cal = 16'b0000010011001011;
            15'd16169: log10_cal = 16'b0000010011001011;
            15'd16170: log10_cal = 16'b0000010011001011;
            15'd16171: log10_cal = 16'b0000010011001011;
            15'd16172: log10_cal = 16'b0000010011001011;
            15'd16173: log10_cal = 16'b0000010011001011;
            15'd16174: log10_cal = 16'b0000010011001011;
            15'd16175: log10_cal = 16'b0000010011001011;
            15'd16176: log10_cal = 16'b0000010011001011;
            15'd16177: log10_cal = 16'b0000010011001011;
            15'd16178: log10_cal = 16'b0000010011001011;
            15'd16179: log10_cal = 16'b0000010011001011;
            15'd16180: log10_cal = 16'b0000010011001011;
            15'd16181: log10_cal = 16'b0000010011001011;
            15'd16182: log10_cal = 16'b0000010011001011;
            15'd16183: log10_cal = 16'b0000010011001011;
            15'd16184: log10_cal = 16'b0000010011001011;
            15'd16185: log10_cal = 16'b0000010011001011;
            15'd16186: log10_cal = 16'b0000010011001011;
            15'd16187: log10_cal = 16'b0000010011001011;
            15'd16188: log10_cal = 16'b0000010011001011;
            15'd16189: log10_cal = 16'b0000010011001011;
            15'd16190: log10_cal = 16'b0000010011001011;
            15'd16191: log10_cal = 16'b0000010011001011;
            15'd16192: log10_cal = 16'b0000010011001011;
            15'd16193: log10_cal = 16'b0000010011001011;
            15'd16194: log10_cal = 16'b0000010011001011;
            15'd16195: log10_cal = 16'b0000010011001011;
            15'd16196: log10_cal = 16'b0000010011001011;
            15'd16197: log10_cal = 16'b0000010011001011;
            15'd16198: log10_cal = 16'b0000010011001011;
            15'd16199: log10_cal = 16'b0000010011001011;
            15'd16200: log10_cal = 16'b0000010011001011;
            15'd16201: log10_cal = 16'b0000010011001100;
            15'd16202: log10_cal = 16'b0000010011001100;
            15'd16203: log10_cal = 16'b0000010011001100;
            15'd16204: log10_cal = 16'b0000010011001100;
            15'd16205: log10_cal = 16'b0000010011001100;
            15'd16206: log10_cal = 16'b0000010011001100;
            15'd16207: log10_cal = 16'b0000010011001100;
            15'd16208: log10_cal = 16'b0000010011001100;
            15'd16209: log10_cal = 16'b0000010011001100;
            15'd16210: log10_cal = 16'b0000010011001100;
            15'd16211: log10_cal = 16'b0000010011001100;
            15'd16212: log10_cal = 16'b0000010011001100;
            15'd16213: log10_cal = 16'b0000010011001100;
            15'd16214: log10_cal = 16'b0000010011001100;
            15'd16215: log10_cal = 16'b0000010011001100;
            15'd16216: log10_cal = 16'b0000010011001100;
            15'd16217: log10_cal = 16'b0000010011001100;
            15'd16218: log10_cal = 16'b0000010011001100;
            15'd16219: log10_cal = 16'b0000010011001100;
            15'd16220: log10_cal = 16'b0000010011001100;
            15'd16221: log10_cal = 16'b0000010011001100;
            15'd16222: log10_cal = 16'b0000010011001100;
            15'd16223: log10_cal = 16'b0000010011001100;
            15'd16224: log10_cal = 16'b0000010011001100;
            15'd16225: log10_cal = 16'b0000010011001100;
            15'd16226: log10_cal = 16'b0000010011001100;
            15'd16227: log10_cal = 16'b0000010011001100;
            15'd16228: log10_cal = 16'b0000010011001100;
            15'd16229: log10_cal = 16'b0000010011001100;
            15'd16230: log10_cal = 16'b0000010011001100;
            15'd16231: log10_cal = 16'b0000010011001100;
            15'd16232: log10_cal = 16'b0000010011001100;
            15'd16233: log10_cal = 16'b0000010011001100;
            15'd16234: log10_cal = 16'b0000010011001100;
            15'd16235: log10_cal = 16'b0000010011001100;
            15'd16236: log10_cal = 16'b0000010011001100;
            15'd16237: log10_cal = 16'b0000010011001101;
            15'd16238: log10_cal = 16'b0000010011001101;
            15'd16239: log10_cal = 16'b0000010011001101;
            15'd16240: log10_cal = 16'b0000010011001101;
            15'd16241: log10_cal = 16'b0000010011001101;
            15'd16242: log10_cal = 16'b0000010011001101;
            15'd16243: log10_cal = 16'b0000010011001101;
            15'd16244: log10_cal = 16'b0000010011001101;
            15'd16245: log10_cal = 16'b0000010011001101;
            15'd16246: log10_cal = 16'b0000010011001101;
            15'd16247: log10_cal = 16'b0000010011001101;
            15'd16248: log10_cal = 16'b0000010011001101;
            15'd16249: log10_cal = 16'b0000010011001101;
            15'd16250: log10_cal = 16'b0000010011001101;
            15'd16251: log10_cal = 16'b0000010011001101;
            15'd16252: log10_cal = 16'b0000010011001101;
            15'd16253: log10_cal = 16'b0000010011001101;
            15'd16254: log10_cal = 16'b0000010011001101;
            15'd16255: log10_cal = 16'b0000010011001101;
            15'd16256: log10_cal = 16'b0000010011001101;
            15'd16257: log10_cal = 16'b0000010011001101;
            15'd16258: log10_cal = 16'b0000010011001101;
            15'd16259: log10_cal = 16'b0000010011001101;
            15'd16260: log10_cal = 16'b0000010011001101;
            15'd16261: log10_cal = 16'b0000010011001101;
            15'd16262: log10_cal = 16'b0000010011001101;
            15'd16263: log10_cal = 16'b0000010011001101;
            15'd16264: log10_cal = 16'b0000010011001101;
            15'd16265: log10_cal = 16'b0000010011001101;
            15'd16266: log10_cal = 16'b0000010011001101;
            15'd16267: log10_cal = 16'b0000010011001101;
            15'd16268: log10_cal = 16'b0000010011001101;
            15'd16269: log10_cal = 16'b0000010011001101;
            15'd16270: log10_cal = 16'b0000010011001101;
            15'd16271: log10_cal = 16'b0000010011001101;
            15'd16272: log10_cal = 16'b0000010011001101;
            15'd16273: log10_cal = 16'b0000010011001101;
            15'd16274: log10_cal = 16'b0000010011001110;
            15'd16275: log10_cal = 16'b0000010011001110;
            15'd16276: log10_cal = 16'b0000010011001110;
            15'd16277: log10_cal = 16'b0000010011001110;
            15'd16278: log10_cal = 16'b0000010011001110;
            15'd16279: log10_cal = 16'b0000010011001110;
            15'd16280: log10_cal = 16'b0000010011001110;
            15'd16281: log10_cal = 16'b0000010011001110;
            15'd16282: log10_cal = 16'b0000010011001110;
            15'd16283: log10_cal = 16'b0000010011001110;
            15'd16284: log10_cal = 16'b0000010011001110;
            15'd16285: log10_cal = 16'b0000010011001110;
            15'd16286: log10_cal = 16'b0000010011001110;
            15'd16287: log10_cal = 16'b0000010011001110;
            15'd16288: log10_cal = 16'b0000010011001110;
            15'd16289: log10_cal = 16'b0000010011001110;
            15'd16290: log10_cal = 16'b0000010011001110;
            15'd16291: log10_cal = 16'b0000010011001110;
            15'd16292: log10_cal = 16'b0000010011001110;
            15'd16293: log10_cal = 16'b0000010011001110;
            15'd16294: log10_cal = 16'b0000010011001110;
            15'd16295: log10_cal = 16'b0000010011001110;
            15'd16296: log10_cal = 16'b0000010011001110;
            15'd16297: log10_cal = 16'b0000010011001110;
            15'd16298: log10_cal = 16'b0000010011001110;
            15'd16299: log10_cal = 16'b0000010011001110;
            15'd16300: log10_cal = 16'b0000010011001110;
            15'd16301: log10_cal = 16'b0000010011001110;
            15'd16302: log10_cal = 16'b0000010011001110;
            15'd16303: log10_cal = 16'b0000010011001110;
            15'd16304: log10_cal = 16'b0000010011001110;
            15'd16305: log10_cal = 16'b0000010011001110;
            15'd16306: log10_cal = 16'b0000010011001110;
            15'd16307: log10_cal = 16'b0000010011001110;
            15'd16308: log10_cal = 16'b0000010011001110;
            15'd16309: log10_cal = 16'b0000010011001110;
            15'd16310: log10_cal = 16'b0000010011001111;
            15'd16311: log10_cal = 16'b0000010011001111;
            15'd16312: log10_cal = 16'b0000010011001111;
            15'd16313: log10_cal = 16'b0000010011001111;
            15'd16314: log10_cal = 16'b0000010011001111;
            15'd16315: log10_cal = 16'b0000010011001111;
            15'd16316: log10_cal = 16'b0000010011001111;
            15'd16317: log10_cal = 16'b0000010011001111;
            15'd16318: log10_cal = 16'b0000010011001111;
            15'd16319: log10_cal = 16'b0000010011001111;
            15'd16320: log10_cal = 16'b0000010011001111;
            15'd16321: log10_cal = 16'b0000010011001111;
            15'd16322: log10_cal = 16'b0000010011001111;
            15'd16323: log10_cal = 16'b0000010011001111;
            15'd16324: log10_cal = 16'b0000010011001111;
            15'd16325: log10_cal = 16'b0000010011001111;
            15'd16326: log10_cal = 16'b0000010011001111;
            15'd16327: log10_cal = 16'b0000010011001111;
            15'd16328: log10_cal = 16'b0000010011001111;
            15'd16329: log10_cal = 16'b0000010011001111;
            15'd16330: log10_cal = 16'b0000010011001111;
            15'd16331: log10_cal = 16'b0000010011001111;
            15'd16332: log10_cal = 16'b0000010011001111;
            15'd16333: log10_cal = 16'b0000010011001111;
            15'd16334: log10_cal = 16'b0000010011001111;
            15'd16335: log10_cal = 16'b0000010011001111;
            15'd16336: log10_cal = 16'b0000010011001111;
            15'd16337: log10_cal = 16'b0000010011001111;
            15'd16338: log10_cal = 16'b0000010011001111;
            15'd16339: log10_cal = 16'b0000010011001111;
            15'd16340: log10_cal = 16'b0000010011001111;
            15'd16341: log10_cal = 16'b0000010011001111;
            15'd16342: log10_cal = 16'b0000010011001111;
            15'd16343: log10_cal = 16'b0000010011001111;
            15'd16344: log10_cal = 16'b0000010011001111;
            15'd16345: log10_cal = 16'b0000010011001111;
            15'd16346: log10_cal = 16'b0000010011001111;
            15'd16347: log10_cal = 16'b0000010011010000;
            15'd16348: log10_cal = 16'b0000010011010000;
            15'd16349: log10_cal = 16'b0000010011010000;
            15'd16350: log10_cal = 16'b0000010011010000;
            15'd16351: log10_cal = 16'b0000010011010000;
            15'd16352: log10_cal = 16'b0000010011010000;
            15'd16353: log10_cal = 16'b0000010011010000;
            15'd16354: log10_cal = 16'b0000010011010000;
            15'd16355: log10_cal = 16'b0000010011010000;
            15'd16356: log10_cal = 16'b0000010011010000;
            15'd16357: log10_cal = 16'b0000010011010000;
            15'd16358: log10_cal = 16'b0000010011010000;
            15'd16359: log10_cal = 16'b0000010011010000;
            15'd16360: log10_cal = 16'b0000010011010000;
            15'd16361: log10_cal = 16'b0000010011010000;
            15'd16362: log10_cal = 16'b0000010011010000;
            15'd16363: log10_cal = 16'b0000010011010000;
            15'd16364: log10_cal = 16'b0000010011010000;
            15'd16365: log10_cal = 16'b0000010011010000;
            15'd16366: log10_cal = 16'b0000010011010000;
            15'd16367: log10_cal = 16'b0000010011010000;
            15'd16368: log10_cal = 16'b0000010011010000;
            15'd16369: log10_cal = 16'b0000010011010000;
            15'd16370: log10_cal = 16'b0000010011010000;
            15'd16371: log10_cal = 16'b0000010011010000;
            15'd16372: log10_cal = 16'b0000010011010000;
            15'd16373: log10_cal = 16'b0000010011010000;
            15'd16374: log10_cal = 16'b0000010011010000;
            15'd16375: log10_cal = 16'b0000010011010000;
            15'd16376: log10_cal = 16'b0000010011010000;
            15'd16377: log10_cal = 16'b0000010011010000;
            15'd16378: log10_cal = 16'b0000010011010000;
            15'd16379: log10_cal = 16'b0000010011010000;
            15'd16380: log10_cal = 16'b0000010011010000;
            15'd16381: log10_cal = 16'b0000010011010000;
            15'd16382: log10_cal = 16'b0000010011010000;
            15'd16383: log10_cal = 16'b0000010011010000;
            15'd16384: log10_cal = 16'b0000010011010001;
            15'd16385: log10_cal = 16'b0000010011010001;
            15'd16386: log10_cal = 16'b0000010011010001;
            15'd16387: log10_cal = 16'b0000010011010001;
            15'd16388: log10_cal = 16'b0000010011010001;
            15'd16389: log10_cal = 16'b0000010011010001;
            15'd16390: log10_cal = 16'b0000010011010001;
            15'd16391: log10_cal = 16'b0000010011010001;
            15'd16392: log10_cal = 16'b0000010011010001;
            15'd16393: log10_cal = 16'b0000010011010001;
            15'd16394: log10_cal = 16'b0000010011010001;
            15'd16395: log10_cal = 16'b0000010011010001;
            15'd16396: log10_cal = 16'b0000010011010001;
            15'd16397: log10_cal = 16'b0000010011010001;
            15'd16398: log10_cal = 16'b0000010011010001;
            15'd16399: log10_cal = 16'b0000010011010001;
            15'd16400: log10_cal = 16'b0000010011010001;
            15'd16401: log10_cal = 16'b0000010011010001;
            15'd16402: log10_cal = 16'b0000010011010001;
            15'd16403: log10_cal = 16'b0000010011010001;
            15'd16404: log10_cal = 16'b0000010011010001;
            15'd16405: log10_cal = 16'b0000010011010001;
            15'd16406: log10_cal = 16'b0000010011010001;
            15'd16407: log10_cal = 16'b0000010011010001;
            15'd16408: log10_cal = 16'b0000010011010001;
            15'd16409: log10_cal = 16'b0000010011010001;
            15'd16410: log10_cal = 16'b0000010011010001;
            15'd16411: log10_cal = 16'b0000010011010001;
            15'd16412: log10_cal = 16'b0000010011010001;
            15'd16413: log10_cal = 16'b0000010011010001;
            15'd16414: log10_cal = 16'b0000010011010001;
            15'd16415: log10_cal = 16'b0000010011010001;
            15'd16416: log10_cal = 16'b0000010011010001;
            15'd16417: log10_cal = 16'b0000010011010001;
            15'd16418: log10_cal = 16'b0000010011010001;
            15'd16419: log10_cal = 16'b0000010011010001;
            15'd16420: log10_cal = 16'b0000010011010001;
            15'd16421: log10_cal = 16'b0000010011010010;
            15'd16422: log10_cal = 16'b0000010011010010;
            15'd16423: log10_cal = 16'b0000010011010010;
            15'd16424: log10_cal = 16'b0000010011010010;
            15'd16425: log10_cal = 16'b0000010011010010;
            15'd16426: log10_cal = 16'b0000010011010010;
            15'd16427: log10_cal = 16'b0000010011010010;
            15'd16428: log10_cal = 16'b0000010011010010;
            15'd16429: log10_cal = 16'b0000010011010010;
            15'd16430: log10_cal = 16'b0000010011010010;
            15'd16431: log10_cal = 16'b0000010011010010;
            15'd16432: log10_cal = 16'b0000010011010010;
            15'd16433: log10_cal = 16'b0000010011010010;
            15'd16434: log10_cal = 16'b0000010011010010;
            15'd16435: log10_cal = 16'b0000010011010010;
            15'd16436: log10_cal = 16'b0000010011010010;
            15'd16437: log10_cal = 16'b0000010011010010;
            15'd16438: log10_cal = 16'b0000010011010010;
            15'd16439: log10_cal = 16'b0000010011010010;
            15'd16440: log10_cal = 16'b0000010011010010;
            15'd16441: log10_cal = 16'b0000010011010010;
            15'd16442: log10_cal = 16'b0000010011010010;
            15'd16443: log10_cal = 16'b0000010011010010;
            15'd16444: log10_cal = 16'b0000010011010010;
            15'd16445: log10_cal = 16'b0000010011010010;
            15'd16446: log10_cal = 16'b0000010011010010;
            15'd16447: log10_cal = 16'b0000010011010010;
            15'd16448: log10_cal = 16'b0000010011010010;
            15'd16449: log10_cal = 16'b0000010011010010;
            15'd16450: log10_cal = 16'b0000010011010010;
            15'd16451: log10_cal = 16'b0000010011010010;
            15'd16452: log10_cal = 16'b0000010011010010;
            15'd16453: log10_cal = 16'b0000010011010010;
            15'd16454: log10_cal = 16'b0000010011010010;
            15'd16455: log10_cal = 16'b0000010011010010;
            15'd16456: log10_cal = 16'b0000010011010010;
            15'd16457: log10_cal = 16'b0000010011010010;
            15'd16458: log10_cal = 16'b0000010011010011;
            15'd16459: log10_cal = 16'b0000010011010011;
            15'd16460: log10_cal = 16'b0000010011010011;
            15'd16461: log10_cal = 16'b0000010011010011;
            15'd16462: log10_cal = 16'b0000010011010011;
            15'd16463: log10_cal = 16'b0000010011010011;
            15'd16464: log10_cal = 16'b0000010011010011;
            15'd16465: log10_cal = 16'b0000010011010011;
            15'd16466: log10_cal = 16'b0000010011010011;
            15'd16467: log10_cal = 16'b0000010011010011;
            15'd16468: log10_cal = 16'b0000010011010011;
            15'd16469: log10_cal = 16'b0000010011010011;
            15'd16470: log10_cal = 16'b0000010011010011;
            15'd16471: log10_cal = 16'b0000010011010011;
            15'd16472: log10_cal = 16'b0000010011010011;
            15'd16473: log10_cal = 16'b0000010011010011;
            15'd16474: log10_cal = 16'b0000010011010011;
            15'd16475: log10_cal = 16'b0000010011010011;
            15'd16476: log10_cal = 16'b0000010011010011;
            15'd16477: log10_cal = 16'b0000010011010011;
            15'd16478: log10_cal = 16'b0000010011010011;
            15'd16479: log10_cal = 16'b0000010011010011;
            15'd16480: log10_cal = 16'b0000010011010011;
            15'd16481: log10_cal = 16'b0000010011010011;
            15'd16482: log10_cal = 16'b0000010011010011;
            15'd16483: log10_cal = 16'b0000010011010011;
            15'd16484: log10_cal = 16'b0000010011010011;
            15'd16485: log10_cal = 16'b0000010011010011;
            15'd16486: log10_cal = 16'b0000010011010011;
            15'd16487: log10_cal = 16'b0000010011010011;
            15'd16488: log10_cal = 16'b0000010011010011;
            15'd16489: log10_cal = 16'b0000010011010011;
            15'd16490: log10_cal = 16'b0000010011010011;
            15'd16491: log10_cal = 16'b0000010011010011;
            15'd16492: log10_cal = 16'b0000010011010011;
            15'd16493: log10_cal = 16'b0000010011010011;
            15'd16494: log10_cal = 16'b0000010011010011;
            15'd16495: log10_cal = 16'b0000010011010100;
            15'd16496: log10_cal = 16'b0000010011010100;
            15'd16497: log10_cal = 16'b0000010011010100;
            15'd16498: log10_cal = 16'b0000010011010100;
            15'd16499: log10_cal = 16'b0000010011010100;
            15'd16500: log10_cal = 16'b0000010011010100;
            15'd16501: log10_cal = 16'b0000010011010100;
            15'd16502: log10_cal = 16'b0000010011010100;
            15'd16503: log10_cal = 16'b0000010011010100;
            15'd16504: log10_cal = 16'b0000010011010100;
            15'd16505: log10_cal = 16'b0000010011010100;
            15'd16506: log10_cal = 16'b0000010011010100;
            15'd16507: log10_cal = 16'b0000010011010100;
            15'd16508: log10_cal = 16'b0000010011010100;
            15'd16509: log10_cal = 16'b0000010011010100;
            15'd16510: log10_cal = 16'b0000010011010100;
            15'd16511: log10_cal = 16'b0000010011010100;
            15'd16512: log10_cal = 16'b0000010011010100;
            15'd16513: log10_cal = 16'b0000010011010100;
            15'd16514: log10_cal = 16'b0000010011010100;
            15'd16515: log10_cal = 16'b0000010011010100;
            15'd16516: log10_cal = 16'b0000010011010100;
            15'd16517: log10_cal = 16'b0000010011010100;
            15'd16518: log10_cal = 16'b0000010011010100;
            15'd16519: log10_cal = 16'b0000010011010100;
            15'd16520: log10_cal = 16'b0000010011010100;
            15'd16521: log10_cal = 16'b0000010011010100;
            15'd16522: log10_cal = 16'b0000010011010100;
            15'd16523: log10_cal = 16'b0000010011010100;
            15'd16524: log10_cal = 16'b0000010011010100;
            15'd16525: log10_cal = 16'b0000010011010100;
            15'd16526: log10_cal = 16'b0000010011010100;
            15'd16527: log10_cal = 16'b0000010011010100;
            15'd16528: log10_cal = 16'b0000010011010100;
            15'd16529: log10_cal = 16'b0000010011010100;
            15'd16530: log10_cal = 16'b0000010011010100;
            15'd16531: log10_cal = 16'b0000010011010100;
            15'd16532: log10_cal = 16'b0000010011010101;
            15'd16533: log10_cal = 16'b0000010011010101;
            15'd16534: log10_cal = 16'b0000010011010101;
            15'd16535: log10_cal = 16'b0000010011010101;
            15'd16536: log10_cal = 16'b0000010011010101;
            15'd16537: log10_cal = 16'b0000010011010101;
            15'd16538: log10_cal = 16'b0000010011010101;
            15'd16539: log10_cal = 16'b0000010011010101;
            15'd16540: log10_cal = 16'b0000010011010101;
            15'd16541: log10_cal = 16'b0000010011010101;
            15'd16542: log10_cal = 16'b0000010011010101;
            15'd16543: log10_cal = 16'b0000010011010101;
            15'd16544: log10_cal = 16'b0000010011010101;
            15'd16545: log10_cal = 16'b0000010011010101;
            15'd16546: log10_cal = 16'b0000010011010101;
            15'd16547: log10_cal = 16'b0000010011010101;
            15'd16548: log10_cal = 16'b0000010011010101;
            15'd16549: log10_cal = 16'b0000010011010101;
            15'd16550: log10_cal = 16'b0000010011010101;
            15'd16551: log10_cal = 16'b0000010011010101;
            15'd16552: log10_cal = 16'b0000010011010101;
            15'd16553: log10_cal = 16'b0000010011010101;
            15'd16554: log10_cal = 16'b0000010011010101;
            15'd16555: log10_cal = 16'b0000010011010101;
            15'd16556: log10_cal = 16'b0000010011010101;
            15'd16557: log10_cal = 16'b0000010011010101;
            15'd16558: log10_cal = 16'b0000010011010101;
            15'd16559: log10_cal = 16'b0000010011010101;
            15'd16560: log10_cal = 16'b0000010011010101;
            15'd16561: log10_cal = 16'b0000010011010101;
            15'd16562: log10_cal = 16'b0000010011010101;
            15'd16563: log10_cal = 16'b0000010011010101;
            15'd16564: log10_cal = 16'b0000010011010101;
            15'd16565: log10_cal = 16'b0000010011010101;
            15'd16566: log10_cal = 16'b0000010011010101;
            15'd16567: log10_cal = 16'b0000010011010101;
            15'd16568: log10_cal = 16'b0000010011010101;
            15'd16569: log10_cal = 16'b0000010011010110;
            15'd16570: log10_cal = 16'b0000010011010110;
            15'd16571: log10_cal = 16'b0000010011010110;
            15'd16572: log10_cal = 16'b0000010011010110;
            15'd16573: log10_cal = 16'b0000010011010110;
            15'd16574: log10_cal = 16'b0000010011010110;
            15'd16575: log10_cal = 16'b0000010011010110;
            15'd16576: log10_cal = 16'b0000010011010110;
            15'd16577: log10_cal = 16'b0000010011010110;
            15'd16578: log10_cal = 16'b0000010011010110;
            15'd16579: log10_cal = 16'b0000010011010110;
            15'd16580: log10_cal = 16'b0000010011010110;
            15'd16581: log10_cal = 16'b0000010011010110;
            15'd16582: log10_cal = 16'b0000010011010110;
            15'd16583: log10_cal = 16'b0000010011010110;
            15'd16584: log10_cal = 16'b0000010011010110;
            15'd16585: log10_cal = 16'b0000010011010110;
            15'd16586: log10_cal = 16'b0000010011010110;
            15'd16587: log10_cal = 16'b0000010011010110;
            15'd16588: log10_cal = 16'b0000010011010110;
            15'd16589: log10_cal = 16'b0000010011010110;
            15'd16590: log10_cal = 16'b0000010011010110;
            15'd16591: log10_cal = 16'b0000010011010110;
            15'd16592: log10_cal = 16'b0000010011010110;
            15'd16593: log10_cal = 16'b0000010011010110;
            15'd16594: log10_cal = 16'b0000010011010110;
            15'd16595: log10_cal = 16'b0000010011010110;
            15'd16596: log10_cal = 16'b0000010011010110;
            15'd16597: log10_cal = 16'b0000010011010110;
            15'd16598: log10_cal = 16'b0000010011010110;
            15'd16599: log10_cal = 16'b0000010011010110;
            15'd16600: log10_cal = 16'b0000010011010110;
            15'd16601: log10_cal = 16'b0000010011010110;
            15'd16602: log10_cal = 16'b0000010011010110;
            15'd16603: log10_cal = 16'b0000010011010110;
            15'd16604: log10_cal = 16'b0000010011010110;
            15'd16605: log10_cal = 16'b0000010011010110;
            15'd16606: log10_cal = 16'b0000010011010111;
            15'd16607: log10_cal = 16'b0000010011010111;
            15'd16608: log10_cal = 16'b0000010011010111;
            15'd16609: log10_cal = 16'b0000010011010111;
            15'd16610: log10_cal = 16'b0000010011010111;
            15'd16611: log10_cal = 16'b0000010011010111;
            15'd16612: log10_cal = 16'b0000010011010111;
            15'd16613: log10_cal = 16'b0000010011010111;
            15'd16614: log10_cal = 16'b0000010011010111;
            15'd16615: log10_cal = 16'b0000010011010111;
            15'd16616: log10_cal = 16'b0000010011010111;
            15'd16617: log10_cal = 16'b0000010011010111;
            15'd16618: log10_cal = 16'b0000010011010111;
            15'd16619: log10_cal = 16'b0000010011010111;
            15'd16620: log10_cal = 16'b0000010011010111;
            15'd16621: log10_cal = 16'b0000010011010111;
            15'd16622: log10_cal = 16'b0000010011010111;
            15'd16623: log10_cal = 16'b0000010011010111;
            15'd16624: log10_cal = 16'b0000010011010111;
            15'd16625: log10_cal = 16'b0000010011010111;
            15'd16626: log10_cal = 16'b0000010011010111;
            15'd16627: log10_cal = 16'b0000010011010111;
            15'd16628: log10_cal = 16'b0000010011010111;
            15'd16629: log10_cal = 16'b0000010011010111;
            15'd16630: log10_cal = 16'b0000010011010111;
            15'd16631: log10_cal = 16'b0000010011010111;
            15'd16632: log10_cal = 16'b0000010011010111;
            15'd16633: log10_cal = 16'b0000010011010111;
            15'd16634: log10_cal = 16'b0000010011010111;
            15'd16635: log10_cal = 16'b0000010011010111;
            15'd16636: log10_cal = 16'b0000010011010111;
            15'd16637: log10_cal = 16'b0000010011010111;
            15'd16638: log10_cal = 16'b0000010011010111;
            15'd16639: log10_cal = 16'b0000010011010111;
            15'd16640: log10_cal = 16'b0000010011010111;
            15'd16641: log10_cal = 16'b0000010011010111;
            15'd16642: log10_cal = 16'b0000010011010111;
            15'd16643: log10_cal = 16'b0000010011010111;
            15'd16644: log10_cal = 16'b0000010011011000;
            15'd16645: log10_cal = 16'b0000010011011000;
            15'd16646: log10_cal = 16'b0000010011011000;
            15'd16647: log10_cal = 16'b0000010011011000;
            15'd16648: log10_cal = 16'b0000010011011000;
            15'd16649: log10_cal = 16'b0000010011011000;
            15'd16650: log10_cal = 16'b0000010011011000;
            15'd16651: log10_cal = 16'b0000010011011000;
            15'd16652: log10_cal = 16'b0000010011011000;
            15'd16653: log10_cal = 16'b0000010011011000;
            15'd16654: log10_cal = 16'b0000010011011000;
            15'd16655: log10_cal = 16'b0000010011011000;
            15'd16656: log10_cal = 16'b0000010011011000;
            15'd16657: log10_cal = 16'b0000010011011000;
            15'd16658: log10_cal = 16'b0000010011011000;
            15'd16659: log10_cal = 16'b0000010011011000;
            15'd16660: log10_cal = 16'b0000010011011000;
            15'd16661: log10_cal = 16'b0000010011011000;
            15'd16662: log10_cal = 16'b0000010011011000;
            15'd16663: log10_cal = 16'b0000010011011000;
            15'd16664: log10_cal = 16'b0000010011011000;
            15'd16665: log10_cal = 16'b0000010011011000;
            15'd16666: log10_cal = 16'b0000010011011000;
            15'd16667: log10_cal = 16'b0000010011011000;
            15'd16668: log10_cal = 16'b0000010011011000;
            15'd16669: log10_cal = 16'b0000010011011000;
            15'd16670: log10_cal = 16'b0000010011011000;
            15'd16671: log10_cal = 16'b0000010011011000;
            15'd16672: log10_cal = 16'b0000010011011000;
            15'd16673: log10_cal = 16'b0000010011011000;
            15'd16674: log10_cal = 16'b0000010011011000;
            15'd16675: log10_cal = 16'b0000010011011000;
            15'd16676: log10_cal = 16'b0000010011011000;
            15'd16677: log10_cal = 16'b0000010011011000;
            15'd16678: log10_cal = 16'b0000010011011000;
            15'd16679: log10_cal = 16'b0000010011011000;
            15'd16680: log10_cal = 16'b0000010011011000;
            15'd16681: log10_cal = 16'b0000010011011001;
            15'd16682: log10_cal = 16'b0000010011011001;
            15'd16683: log10_cal = 16'b0000010011011001;
            15'd16684: log10_cal = 16'b0000010011011001;
            15'd16685: log10_cal = 16'b0000010011011001;
            15'd16686: log10_cal = 16'b0000010011011001;
            15'd16687: log10_cal = 16'b0000010011011001;
            15'd16688: log10_cal = 16'b0000010011011001;
            15'd16689: log10_cal = 16'b0000010011011001;
            15'd16690: log10_cal = 16'b0000010011011001;
            15'd16691: log10_cal = 16'b0000010011011001;
            15'd16692: log10_cal = 16'b0000010011011001;
            15'd16693: log10_cal = 16'b0000010011011001;
            15'd16694: log10_cal = 16'b0000010011011001;
            15'd16695: log10_cal = 16'b0000010011011001;
            15'd16696: log10_cal = 16'b0000010011011001;
            15'd16697: log10_cal = 16'b0000010011011001;
            15'd16698: log10_cal = 16'b0000010011011001;
            15'd16699: log10_cal = 16'b0000010011011001;
            15'd16700: log10_cal = 16'b0000010011011001;
            15'd16701: log10_cal = 16'b0000010011011001;
            15'd16702: log10_cal = 16'b0000010011011001;
            15'd16703: log10_cal = 16'b0000010011011001;
            15'd16704: log10_cal = 16'b0000010011011001;
            15'd16705: log10_cal = 16'b0000010011011001;
            15'd16706: log10_cal = 16'b0000010011011001;
            15'd16707: log10_cal = 16'b0000010011011001;
            15'd16708: log10_cal = 16'b0000010011011001;
            15'd16709: log10_cal = 16'b0000010011011001;
            15'd16710: log10_cal = 16'b0000010011011001;
            15'd16711: log10_cal = 16'b0000010011011001;
            15'd16712: log10_cal = 16'b0000010011011001;
            15'd16713: log10_cal = 16'b0000010011011001;
            15'd16714: log10_cal = 16'b0000010011011001;
            15'd16715: log10_cal = 16'b0000010011011001;
            15'd16716: log10_cal = 16'b0000010011011001;
            15'd16717: log10_cal = 16'b0000010011011001;
            15'd16718: log10_cal = 16'b0000010011011001;
            15'd16719: log10_cal = 16'b0000010011011010;
            15'd16720: log10_cal = 16'b0000010011011010;
            15'd16721: log10_cal = 16'b0000010011011010;
            15'd16722: log10_cal = 16'b0000010011011010;
            15'd16723: log10_cal = 16'b0000010011011010;
            15'd16724: log10_cal = 16'b0000010011011010;
            15'd16725: log10_cal = 16'b0000010011011010;
            15'd16726: log10_cal = 16'b0000010011011010;
            15'd16727: log10_cal = 16'b0000010011011010;
            15'd16728: log10_cal = 16'b0000010011011010;
            15'd16729: log10_cal = 16'b0000010011011010;
            15'd16730: log10_cal = 16'b0000010011011010;
            15'd16731: log10_cal = 16'b0000010011011010;
            15'd16732: log10_cal = 16'b0000010011011010;
            15'd16733: log10_cal = 16'b0000010011011010;
            15'd16734: log10_cal = 16'b0000010011011010;
            15'd16735: log10_cal = 16'b0000010011011010;
            15'd16736: log10_cal = 16'b0000010011011010;
            15'd16737: log10_cal = 16'b0000010011011010;
            15'd16738: log10_cal = 16'b0000010011011010;
            15'd16739: log10_cal = 16'b0000010011011010;
            15'd16740: log10_cal = 16'b0000010011011010;
            15'd16741: log10_cal = 16'b0000010011011010;
            15'd16742: log10_cal = 16'b0000010011011010;
            15'd16743: log10_cal = 16'b0000010011011010;
            15'd16744: log10_cal = 16'b0000010011011010;
            15'd16745: log10_cal = 16'b0000010011011010;
            15'd16746: log10_cal = 16'b0000010011011010;
            15'd16747: log10_cal = 16'b0000010011011010;
            15'd16748: log10_cal = 16'b0000010011011010;
            15'd16749: log10_cal = 16'b0000010011011010;
            15'd16750: log10_cal = 16'b0000010011011010;
            15'd16751: log10_cal = 16'b0000010011011010;
            15'd16752: log10_cal = 16'b0000010011011010;
            15'd16753: log10_cal = 16'b0000010011011010;
            15'd16754: log10_cal = 16'b0000010011011010;
            15'd16755: log10_cal = 16'b0000010011011010;
            15'd16756: log10_cal = 16'b0000010011011011;
            15'd16757: log10_cal = 16'b0000010011011011;
            15'd16758: log10_cal = 16'b0000010011011011;
            15'd16759: log10_cal = 16'b0000010011011011;
            15'd16760: log10_cal = 16'b0000010011011011;
            15'd16761: log10_cal = 16'b0000010011011011;
            15'd16762: log10_cal = 16'b0000010011011011;
            15'd16763: log10_cal = 16'b0000010011011011;
            15'd16764: log10_cal = 16'b0000010011011011;
            15'd16765: log10_cal = 16'b0000010011011011;
            15'd16766: log10_cal = 16'b0000010011011011;
            15'd16767: log10_cal = 16'b0000010011011011;
            15'd16768: log10_cal = 16'b0000010011011011;
            15'd16769: log10_cal = 16'b0000010011011011;
            15'd16770: log10_cal = 16'b0000010011011011;
            15'd16771: log10_cal = 16'b0000010011011011;
            15'd16772: log10_cal = 16'b0000010011011011;
            15'd16773: log10_cal = 16'b0000010011011011;
            15'd16774: log10_cal = 16'b0000010011011011;
            15'd16775: log10_cal = 16'b0000010011011011;
            15'd16776: log10_cal = 16'b0000010011011011;
            15'd16777: log10_cal = 16'b0000010011011011;
            15'd16778: log10_cal = 16'b0000010011011011;
            15'd16779: log10_cal = 16'b0000010011011011;
            15'd16780: log10_cal = 16'b0000010011011011;
            15'd16781: log10_cal = 16'b0000010011011011;
            15'd16782: log10_cal = 16'b0000010011011011;
            15'd16783: log10_cal = 16'b0000010011011011;
            15'd16784: log10_cal = 16'b0000010011011011;
            15'd16785: log10_cal = 16'b0000010011011011;
            15'd16786: log10_cal = 16'b0000010011011011;
            15'd16787: log10_cal = 16'b0000010011011011;
            15'd16788: log10_cal = 16'b0000010011011011;
            15'd16789: log10_cal = 16'b0000010011011011;
            15'd16790: log10_cal = 16'b0000010011011011;
            15'd16791: log10_cal = 16'b0000010011011011;
            15'd16792: log10_cal = 16'b0000010011011011;
            15'd16793: log10_cal = 16'b0000010011011011;
            15'd16794: log10_cal = 16'b0000010011011100;
            15'd16795: log10_cal = 16'b0000010011011100;
            15'd16796: log10_cal = 16'b0000010011011100;
            15'd16797: log10_cal = 16'b0000010011011100;
            15'd16798: log10_cal = 16'b0000010011011100;
            15'd16799: log10_cal = 16'b0000010011011100;
            15'd16800: log10_cal = 16'b0000010011011100;
            15'd16801: log10_cal = 16'b0000010011011100;
            15'd16802: log10_cal = 16'b0000010011011100;
            15'd16803: log10_cal = 16'b0000010011011100;
            15'd16804: log10_cal = 16'b0000010011011100;
            15'd16805: log10_cal = 16'b0000010011011100;
            15'd16806: log10_cal = 16'b0000010011011100;
            15'd16807: log10_cal = 16'b0000010011011100;
            15'd16808: log10_cal = 16'b0000010011011100;
            15'd16809: log10_cal = 16'b0000010011011100;
            15'd16810: log10_cal = 16'b0000010011011100;
            15'd16811: log10_cal = 16'b0000010011011100;
            15'd16812: log10_cal = 16'b0000010011011100;
            15'd16813: log10_cal = 16'b0000010011011100;
            15'd16814: log10_cal = 16'b0000010011011100;
            15'd16815: log10_cal = 16'b0000010011011100;
            15'd16816: log10_cal = 16'b0000010011011100;
            15'd16817: log10_cal = 16'b0000010011011100;
            15'd16818: log10_cal = 16'b0000010011011100;
            15'd16819: log10_cal = 16'b0000010011011100;
            15'd16820: log10_cal = 16'b0000010011011100;
            15'd16821: log10_cal = 16'b0000010011011100;
            15'd16822: log10_cal = 16'b0000010011011100;
            15'd16823: log10_cal = 16'b0000010011011100;
            15'd16824: log10_cal = 16'b0000010011011100;
            15'd16825: log10_cal = 16'b0000010011011100;
            15'd16826: log10_cal = 16'b0000010011011100;
            15'd16827: log10_cal = 16'b0000010011011100;
            15'd16828: log10_cal = 16'b0000010011011100;
            15'd16829: log10_cal = 16'b0000010011011100;
            15'd16830: log10_cal = 16'b0000010011011100;
            15'd16831: log10_cal = 16'b0000010011011100;
            15'd16832: log10_cal = 16'b0000010011011101;
            15'd16833: log10_cal = 16'b0000010011011101;
            15'd16834: log10_cal = 16'b0000010011011101;
            15'd16835: log10_cal = 16'b0000010011011101;
            15'd16836: log10_cal = 16'b0000010011011101;
            15'd16837: log10_cal = 16'b0000010011011101;
            15'd16838: log10_cal = 16'b0000010011011101;
            15'd16839: log10_cal = 16'b0000010011011101;
            15'd16840: log10_cal = 16'b0000010011011101;
            15'd16841: log10_cal = 16'b0000010011011101;
            15'd16842: log10_cal = 16'b0000010011011101;
            15'd16843: log10_cal = 16'b0000010011011101;
            15'd16844: log10_cal = 16'b0000010011011101;
            15'd16845: log10_cal = 16'b0000010011011101;
            15'd16846: log10_cal = 16'b0000010011011101;
            15'd16847: log10_cal = 16'b0000010011011101;
            15'd16848: log10_cal = 16'b0000010011011101;
            15'd16849: log10_cal = 16'b0000010011011101;
            15'd16850: log10_cal = 16'b0000010011011101;
            15'd16851: log10_cal = 16'b0000010011011101;
            15'd16852: log10_cal = 16'b0000010011011101;
            15'd16853: log10_cal = 16'b0000010011011101;
            15'd16854: log10_cal = 16'b0000010011011101;
            15'd16855: log10_cal = 16'b0000010011011101;
            15'd16856: log10_cal = 16'b0000010011011101;
            15'd16857: log10_cal = 16'b0000010011011101;
            15'd16858: log10_cal = 16'b0000010011011101;
            15'd16859: log10_cal = 16'b0000010011011101;
            15'd16860: log10_cal = 16'b0000010011011101;
            15'd16861: log10_cal = 16'b0000010011011101;
            15'd16862: log10_cal = 16'b0000010011011101;
            15'd16863: log10_cal = 16'b0000010011011101;
            15'd16864: log10_cal = 16'b0000010011011101;
            15'd16865: log10_cal = 16'b0000010011011101;
            15'd16866: log10_cal = 16'b0000010011011101;
            15'd16867: log10_cal = 16'b0000010011011101;
            15'd16868: log10_cal = 16'b0000010011011101;
            15'd16869: log10_cal = 16'b0000010011011101;
            15'd16870: log10_cal = 16'b0000010011011110;
            15'd16871: log10_cal = 16'b0000010011011110;
            15'd16872: log10_cal = 16'b0000010011011110;
            15'd16873: log10_cal = 16'b0000010011011110;
            15'd16874: log10_cal = 16'b0000010011011110;
            15'd16875: log10_cal = 16'b0000010011011110;
            15'd16876: log10_cal = 16'b0000010011011110;
            15'd16877: log10_cal = 16'b0000010011011110;
            15'd16878: log10_cal = 16'b0000010011011110;
            15'd16879: log10_cal = 16'b0000010011011110;
            15'd16880: log10_cal = 16'b0000010011011110;
            15'd16881: log10_cal = 16'b0000010011011110;
            15'd16882: log10_cal = 16'b0000010011011110;
            15'd16883: log10_cal = 16'b0000010011011110;
            15'd16884: log10_cal = 16'b0000010011011110;
            15'd16885: log10_cal = 16'b0000010011011110;
            15'd16886: log10_cal = 16'b0000010011011110;
            15'd16887: log10_cal = 16'b0000010011011110;
            15'd16888: log10_cal = 16'b0000010011011110;
            15'd16889: log10_cal = 16'b0000010011011110;
            15'd16890: log10_cal = 16'b0000010011011110;
            15'd16891: log10_cal = 16'b0000010011011110;
            15'd16892: log10_cal = 16'b0000010011011110;
            15'd16893: log10_cal = 16'b0000010011011110;
            15'd16894: log10_cal = 16'b0000010011011110;
            15'd16895: log10_cal = 16'b0000010011011110;
            15'd16896: log10_cal = 16'b0000010011011110;
            15'd16897: log10_cal = 16'b0000010011011110;
            15'd16898: log10_cal = 16'b0000010011011110;
            15'd16899: log10_cal = 16'b0000010011011110;
            15'd16900: log10_cal = 16'b0000010011011110;
            15'd16901: log10_cal = 16'b0000010011011110;
            15'd16902: log10_cal = 16'b0000010011011110;
            15'd16903: log10_cal = 16'b0000010011011110;
            15'd16904: log10_cal = 16'b0000010011011110;
            15'd16905: log10_cal = 16'b0000010011011110;
            15'd16906: log10_cal = 16'b0000010011011110;
            15'd16907: log10_cal = 16'b0000010011011110;
            15'd16908: log10_cal = 16'b0000010011011111;
            15'd16909: log10_cal = 16'b0000010011011111;
            15'd16910: log10_cal = 16'b0000010011011111;
            15'd16911: log10_cal = 16'b0000010011011111;
            15'd16912: log10_cal = 16'b0000010011011111;
            15'd16913: log10_cal = 16'b0000010011011111;
            15'd16914: log10_cal = 16'b0000010011011111;
            15'd16915: log10_cal = 16'b0000010011011111;
            15'd16916: log10_cal = 16'b0000010011011111;
            15'd16917: log10_cal = 16'b0000010011011111;
            15'd16918: log10_cal = 16'b0000010011011111;
            15'd16919: log10_cal = 16'b0000010011011111;
            15'd16920: log10_cal = 16'b0000010011011111;
            15'd16921: log10_cal = 16'b0000010011011111;
            15'd16922: log10_cal = 16'b0000010011011111;
            15'd16923: log10_cal = 16'b0000010011011111;
            15'd16924: log10_cal = 16'b0000010011011111;
            15'd16925: log10_cal = 16'b0000010011011111;
            15'd16926: log10_cal = 16'b0000010011011111;
            15'd16927: log10_cal = 16'b0000010011011111;
            15'd16928: log10_cal = 16'b0000010011011111;
            15'd16929: log10_cal = 16'b0000010011011111;
            15'd16930: log10_cal = 16'b0000010011011111;
            15'd16931: log10_cal = 16'b0000010011011111;
            15'd16932: log10_cal = 16'b0000010011011111;
            15'd16933: log10_cal = 16'b0000010011011111;
            15'd16934: log10_cal = 16'b0000010011011111;
            15'd16935: log10_cal = 16'b0000010011011111;
            15'd16936: log10_cal = 16'b0000010011011111;
            15'd16937: log10_cal = 16'b0000010011011111;
            15'd16938: log10_cal = 16'b0000010011011111;
            15'd16939: log10_cal = 16'b0000010011011111;
            15'd16940: log10_cal = 16'b0000010011011111;
            15'd16941: log10_cal = 16'b0000010011011111;
            15'd16942: log10_cal = 16'b0000010011011111;
            15'd16943: log10_cal = 16'b0000010011011111;
            15'd16944: log10_cal = 16'b0000010011011111;
            15'd16945: log10_cal = 16'b0000010011011111;
            15'd16946: log10_cal = 16'b0000010011100000;
            15'd16947: log10_cal = 16'b0000010011100000;
            15'd16948: log10_cal = 16'b0000010011100000;
            15'd16949: log10_cal = 16'b0000010011100000;
            15'd16950: log10_cal = 16'b0000010011100000;
            15'd16951: log10_cal = 16'b0000010011100000;
            15'd16952: log10_cal = 16'b0000010011100000;
            15'd16953: log10_cal = 16'b0000010011100000;
            15'd16954: log10_cal = 16'b0000010011100000;
            15'd16955: log10_cal = 16'b0000010011100000;
            15'd16956: log10_cal = 16'b0000010011100000;
            15'd16957: log10_cal = 16'b0000010011100000;
            15'd16958: log10_cal = 16'b0000010011100000;
            15'd16959: log10_cal = 16'b0000010011100000;
            15'd16960: log10_cal = 16'b0000010011100000;
            15'd16961: log10_cal = 16'b0000010011100000;
            15'd16962: log10_cal = 16'b0000010011100000;
            15'd16963: log10_cal = 16'b0000010011100000;
            15'd16964: log10_cal = 16'b0000010011100000;
            15'd16965: log10_cal = 16'b0000010011100000;
            15'd16966: log10_cal = 16'b0000010011100000;
            15'd16967: log10_cal = 16'b0000010011100000;
            15'd16968: log10_cal = 16'b0000010011100000;
            15'd16969: log10_cal = 16'b0000010011100000;
            15'd16970: log10_cal = 16'b0000010011100000;
            15'd16971: log10_cal = 16'b0000010011100000;
            15'd16972: log10_cal = 16'b0000010011100000;
            15'd16973: log10_cal = 16'b0000010011100000;
            15'd16974: log10_cal = 16'b0000010011100000;
            15'd16975: log10_cal = 16'b0000010011100000;
            15'd16976: log10_cal = 16'b0000010011100000;
            15'd16977: log10_cal = 16'b0000010011100000;
            15'd16978: log10_cal = 16'b0000010011100000;
            15'd16979: log10_cal = 16'b0000010011100000;
            15'd16980: log10_cal = 16'b0000010011100000;
            15'd16981: log10_cal = 16'b0000010011100000;
            15'd16982: log10_cal = 16'b0000010011100000;
            15'd16983: log10_cal = 16'b0000010011100000;
            15'd16984: log10_cal = 16'b0000010011100001;
            15'd16985: log10_cal = 16'b0000010011100001;
            15'd16986: log10_cal = 16'b0000010011100001;
            15'd16987: log10_cal = 16'b0000010011100001;
            15'd16988: log10_cal = 16'b0000010011100001;
            15'd16989: log10_cal = 16'b0000010011100001;
            15'd16990: log10_cal = 16'b0000010011100001;
            15'd16991: log10_cal = 16'b0000010011100001;
            15'd16992: log10_cal = 16'b0000010011100001;
            15'd16993: log10_cal = 16'b0000010011100001;
            15'd16994: log10_cal = 16'b0000010011100001;
            15'd16995: log10_cal = 16'b0000010011100001;
            15'd16996: log10_cal = 16'b0000010011100001;
            15'd16997: log10_cal = 16'b0000010011100001;
            15'd16998: log10_cal = 16'b0000010011100001;
            15'd16999: log10_cal = 16'b0000010011100001;
            15'd17000: log10_cal = 16'b0000010011100001;
            15'd17001: log10_cal = 16'b0000010011100001;
            15'd17002: log10_cal = 16'b0000010011100001;
            15'd17003: log10_cal = 16'b0000010011100001;
            15'd17004: log10_cal = 16'b0000010011100001;
            15'd17005: log10_cal = 16'b0000010011100001;
            15'd17006: log10_cal = 16'b0000010011100001;
            15'd17007: log10_cal = 16'b0000010011100001;
            15'd17008: log10_cal = 16'b0000010011100001;
            15'd17009: log10_cal = 16'b0000010011100001;
            15'd17010: log10_cal = 16'b0000010011100001;
            15'd17011: log10_cal = 16'b0000010011100001;
            15'd17012: log10_cal = 16'b0000010011100001;
            15'd17013: log10_cal = 16'b0000010011100001;
            15'd17014: log10_cal = 16'b0000010011100001;
            15'd17015: log10_cal = 16'b0000010011100001;
            15'd17016: log10_cal = 16'b0000010011100001;
            15'd17017: log10_cal = 16'b0000010011100001;
            15'd17018: log10_cal = 16'b0000010011100001;
            15'd17019: log10_cal = 16'b0000010011100001;
            15'd17020: log10_cal = 16'b0000010011100001;
            15'd17021: log10_cal = 16'b0000010011100001;
            15'd17022: log10_cal = 16'b0000010011100010;
            15'd17023: log10_cal = 16'b0000010011100010;
            15'd17024: log10_cal = 16'b0000010011100010;
            15'd17025: log10_cal = 16'b0000010011100010;
            15'd17026: log10_cal = 16'b0000010011100010;
            15'd17027: log10_cal = 16'b0000010011100010;
            15'd17028: log10_cal = 16'b0000010011100010;
            15'd17029: log10_cal = 16'b0000010011100010;
            15'd17030: log10_cal = 16'b0000010011100010;
            15'd17031: log10_cal = 16'b0000010011100010;
            15'd17032: log10_cal = 16'b0000010011100010;
            15'd17033: log10_cal = 16'b0000010011100010;
            15'd17034: log10_cal = 16'b0000010011100010;
            15'd17035: log10_cal = 16'b0000010011100010;
            15'd17036: log10_cal = 16'b0000010011100010;
            15'd17037: log10_cal = 16'b0000010011100010;
            15'd17038: log10_cal = 16'b0000010011100010;
            15'd17039: log10_cal = 16'b0000010011100010;
            15'd17040: log10_cal = 16'b0000010011100010;
            15'd17041: log10_cal = 16'b0000010011100010;
            15'd17042: log10_cal = 16'b0000010011100010;
            15'd17043: log10_cal = 16'b0000010011100010;
            15'd17044: log10_cal = 16'b0000010011100010;
            15'd17045: log10_cal = 16'b0000010011100010;
            15'd17046: log10_cal = 16'b0000010011100010;
            15'd17047: log10_cal = 16'b0000010011100010;
            15'd17048: log10_cal = 16'b0000010011100010;
            15'd17049: log10_cal = 16'b0000010011100010;
            15'd17050: log10_cal = 16'b0000010011100010;
            15'd17051: log10_cal = 16'b0000010011100010;
            15'd17052: log10_cal = 16'b0000010011100010;
            15'd17053: log10_cal = 16'b0000010011100010;
            15'd17054: log10_cal = 16'b0000010011100010;
            15'd17055: log10_cal = 16'b0000010011100010;
            15'd17056: log10_cal = 16'b0000010011100010;
            15'd17057: log10_cal = 16'b0000010011100010;
            15'd17058: log10_cal = 16'b0000010011100010;
            15'd17059: log10_cal = 16'b0000010011100010;
            15'd17060: log10_cal = 16'b0000010011100010;
            15'd17061: log10_cal = 16'b0000010011100011;
            15'd17062: log10_cal = 16'b0000010011100011;
            15'd17063: log10_cal = 16'b0000010011100011;
            15'd17064: log10_cal = 16'b0000010011100011;
            15'd17065: log10_cal = 16'b0000010011100011;
            15'd17066: log10_cal = 16'b0000010011100011;
            15'd17067: log10_cal = 16'b0000010011100011;
            15'd17068: log10_cal = 16'b0000010011100011;
            15'd17069: log10_cal = 16'b0000010011100011;
            15'd17070: log10_cal = 16'b0000010011100011;
            15'd17071: log10_cal = 16'b0000010011100011;
            15'd17072: log10_cal = 16'b0000010011100011;
            15'd17073: log10_cal = 16'b0000010011100011;
            15'd17074: log10_cal = 16'b0000010011100011;
            15'd17075: log10_cal = 16'b0000010011100011;
            15'd17076: log10_cal = 16'b0000010011100011;
            15'd17077: log10_cal = 16'b0000010011100011;
            15'd17078: log10_cal = 16'b0000010011100011;
            15'd17079: log10_cal = 16'b0000010011100011;
            15'd17080: log10_cal = 16'b0000010011100011;
            15'd17081: log10_cal = 16'b0000010011100011;
            15'd17082: log10_cal = 16'b0000010011100011;
            15'd17083: log10_cal = 16'b0000010011100011;
            15'd17084: log10_cal = 16'b0000010011100011;
            15'd17085: log10_cal = 16'b0000010011100011;
            15'd17086: log10_cal = 16'b0000010011100011;
            15'd17087: log10_cal = 16'b0000010011100011;
            15'd17088: log10_cal = 16'b0000010011100011;
            15'd17089: log10_cal = 16'b0000010011100011;
            15'd17090: log10_cal = 16'b0000010011100011;
            15'd17091: log10_cal = 16'b0000010011100011;
            15'd17092: log10_cal = 16'b0000010011100011;
            15'd17093: log10_cal = 16'b0000010011100011;
            15'd17094: log10_cal = 16'b0000010011100011;
            15'd17095: log10_cal = 16'b0000010011100011;
            15'd17096: log10_cal = 16'b0000010011100011;
            15'd17097: log10_cal = 16'b0000010011100011;
            15'd17098: log10_cal = 16'b0000010011100011;
            15'd17099: log10_cal = 16'b0000010011100100;
            15'd17100: log10_cal = 16'b0000010011100100;
            15'd17101: log10_cal = 16'b0000010011100100;
            15'd17102: log10_cal = 16'b0000010011100100;
            15'd17103: log10_cal = 16'b0000010011100100;
            15'd17104: log10_cal = 16'b0000010011100100;
            15'd17105: log10_cal = 16'b0000010011100100;
            15'd17106: log10_cal = 16'b0000010011100100;
            15'd17107: log10_cal = 16'b0000010011100100;
            15'd17108: log10_cal = 16'b0000010011100100;
            15'd17109: log10_cal = 16'b0000010011100100;
            15'd17110: log10_cal = 16'b0000010011100100;
            15'd17111: log10_cal = 16'b0000010011100100;
            15'd17112: log10_cal = 16'b0000010011100100;
            15'd17113: log10_cal = 16'b0000010011100100;
            15'd17114: log10_cal = 16'b0000010011100100;
            15'd17115: log10_cal = 16'b0000010011100100;
            15'd17116: log10_cal = 16'b0000010011100100;
            15'd17117: log10_cal = 16'b0000010011100100;
            15'd17118: log10_cal = 16'b0000010011100100;
            15'd17119: log10_cal = 16'b0000010011100100;
            15'd17120: log10_cal = 16'b0000010011100100;
            15'd17121: log10_cal = 16'b0000010011100100;
            15'd17122: log10_cal = 16'b0000010011100100;
            15'd17123: log10_cal = 16'b0000010011100100;
            15'd17124: log10_cal = 16'b0000010011100100;
            15'd17125: log10_cal = 16'b0000010011100100;
            15'd17126: log10_cal = 16'b0000010011100100;
            15'd17127: log10_cal = 16'b0000010011100100;
            15'd17128: log10_cal = 16'b0000010011100100;
            15'd17129: log10_cal = 16'b0000010011100100;
            15'd17130: log10_cal = 16'b0000010011100100;
            15'd17131: log10_cal = 16'b0000010011100100;
            15'd17132: log10_cal = 16'b0000010011100100;
            15'd17133: log10_cal = 16'b0000010011100100;
            15'd17134: log10_cal = 16'b0000010011100100;
            15'd17135: log10_cal = 16'b0000010011100100;
            15'd17136: log10_cal = 16'b0000010011100100;
            15'd17137: log10_cal = 16'b0000010011100101;
            15'd17138: log10_cal = 16'b0000010011100101;
            15'd17139: log10_cal = 16'b0000010011100101;
            15'd17140: log10_cal = 16'b0000010011100101;
            15'd17141: log10_cal = 16'b0000010011100101;
            15'd17142: log10_cal = 16'b0000010011100101;
            15'd17143: log10_cal = 16'b0000010011100101;
            15'd17144: log10_cal = 16'b0000010011100101;
            15'd17145: log10_cal = 16'b0000010011100101;
            15'd17146: log10_cal = 16'b0000010011100101;
            15'd17147: log10_cal = 16'b0000010011100101;
            15'd17148: log10_cal = 16'b0000010011100101;
            15'd17149: log10_cal = 16'b0000010011100101;
            15'd17150: log10_cal = 16'b0000010011100101;
            15'd17151: log10_cal = 16'b0000010011100101;
            15'd17152: log10_cal = 16'b0000010011100101;
            15'd17153: log10_cal = 16'b0000010011100101;
            15'd17154: log10_cal = 16'b0000010011100101;
            15'd17155: log10_cal = 16'b0000010011100101;
            15'd17156: log10_cal = 16'b0000010011100101;
            15'd17157: log10_cal = 16'b0000010011100101;
            15'd17158: log10_cal = 16'b0000010011100101;
            15'd17159: log10_cal = 16'b0000010011100101;
            15'd17160: log10_cal = 16'b0000010011100101;
            15'd17161: log10_cal = 16'b0000010011100101;
            15'd17162: log10_cal = 16'b0000010011100101;
            15'd17163: log10_cal = 16'b0000010011100101;
            15'd17164: log10_cal = 16'b0000010011100101;
            15'd17165: log10_cal = 16'b0000010011100101;
            15'd17166: log10_cal = 16'b0000010011100101;
            15'd17167: log10_cal = 16'b0000010011100101;
            15'd17168: log10_cal = 16'b0000010011100101;
            15'd17169: log10_cal = 16'b0000010011100101;
            15'd17170: log10_cal = 16'b0000010011100101;
            15'd17171: log10_cal = 16'b0000010011100101;
            15'd17172: log10_cal = 16'b0000010011100101;
            15'd17173: log10_cal = 16'b0000010011100101;
            15'd17174: log10_cal = 16'b0000010011100101;
            15'd17175: log10_cal = 16'b0000010011100101;
            15'd17176: log10_cal = 16'b0000010011100110;
            15'd17177: log10_cal = 16'b0000010011100110;
            15'd17178: log10_cal = 16'b0000010011100110;
            15'd17179: log10_cal = 16'b0000010011100110;
            15'd17180: log10_cal = 16'b0000010011100110;
            15'd17181: log10_cal = 16'b0000010011100110;
            15'd17182: log10_cal = 16'b0000010011100110;
            15'd17183: log10_cal = 16'b0000010011100110;
            15'd17184: log10_cal = 16'b0000010011100110;
            15'd17185: log10_cal = 16'b0000010011100110;
            15'd17186: log10_cal = 16'b0000010011100110;
            15'd17187: log10_cal = 16'b0000010011100110;
            15'd17188: log10_cal = 16'b0000010011100110;
            15'd17189: log10_cal = 16'b0000010011100110;
            15'd17190: log10_cal = 16'b0000010011100110;
            15'd17191: log10_cal = 16'b0000010011100110;
            15'd17192: log10_cal = 16'b0000010011100110;
            15'd17193: log10_cal = 16'b0000010011100110;
            15'd17194: log10_cal = 16'b0000010011100110;
            15'd17195: log10_cal = 16'b0000010011100110;
            15'd17196: log10_cal = 16'b0000010011100110;
            15'd17197: log10_cal = 16'b0000010011100110;
            15'd17198: log10_cal = 16'b0000010011100110;
            15'd17199: log10_cal = 16'b0000010011100110;
            15'd17200: log10_cal = 16'b0000010011100110;
            15'd17201: log10_cal = 16'b0000010011100110;
            15'd17202: log10_cal = 16'b0000010011100110;
            15'd17203: log10_cal = 16'b0000010011100110;
            15'd17204: log10_cal = 16'b0000010011100110;
            15'd17205: log10_cal = 16'b0000010011100110;
            15'd17206: log10_cal = 16'b0000010011100110;
            15'd17207: log10_cal = 16'b0000010011100110;
            15'd17208: log10_cal = 16'b0000010011100110;
            15'd17209: log10_cal = 16'b0000010011100110;
            15'd17210: log10_cal = 16'b0000010011100110;
            15'd17211: log10_cal = 16'b0000010011100110;
            15'd17212: log10_cal = 16'b0000010011100110;
            15'd17213: log10_cal = 16'b0000010011100110;
            15'd17214: log10_cal = 16'b0000010011100110;
            15'd17215: log10_cal = 16'b0000010011100111;
            15'd17216: log10_cal = 16'b0000010011100111;
            15'd17217: log10_cal = 16'b0000010011100111;
            15'd17218: log10_cal = 16'b0000010011100111;
            15'd17219: log10_cal = 16'b0000010011100111;
            15'd17220: log10_cal = 16'b0000010011100111;
            15'd17221: log10_cal = 16'b0000010011100111;
            15'd17222: log10_cal = 16'b0000010011100111;
            15'd17223: log10_cal = 16'b0000010011100111;
            15'd17224: log10_cal = 16'b0000010011100111;
            15'd17225: log10_cal = 16'b0000010011100111;
            15'd17226: log10_cal = 16'b0000010011100111;
            15'd17227: log10_cal = 16'b0000010011100111;
            15'd17228: log10_cal = 16'b0000010011100111;
            15'd17229: log10_cal = 16'b0000010011100111;
            15'd17230: log10_cal = 16'b0000010011100111;
            15'd17231: log10_cal = 16'b0000010011100111;
            15'd17232: log10_cal = 16'b0000010011100111;
            15'd17233: log10_cal = 16'b0000010011100111;
            15'd17234: log10_cal = 16'b0000010011100111;
            15'd17235: log10_cal = 16'b0000010011100111;
            15'd17236: log10_cal = 16'b0000010011100111;
            15'd17237: log10_cal = 16'b0000010011100111;
            15'd17238: log10_cal = 16'b0000010011100111;
            15'd17239: log10_cal = 16'b0000010011100111;
            15'd17240: log10_cal = 16'b0000010011100111;
            15'd17241: log10_cal = 16'b0000010011100111;
            15'd17242: log10_cal = 16'b0000010011100111;
            15'd17243: log10_cal = 16'b0000010011100111;
            15'd17244: log10_cal = 16'b0000010011100111;
            15'd17245: log10_cal = 16'b0000010011100111;
            15'd17246: log10_cal = 16'b0000010011100111;
            15'd17247: log10_cal = 16'b0000010011100111;
            15'd17248: log10_cal = 16'b0000010011100111;
            15'd17249: log10_cal = 16'b0000010011100111;
            15'd17250: log10_cal = 16'b0000010011100111;
            15'd17251: log10_cal = 16'b0000010011100111;
            15'd17252: log10_cal = 16'b0000010011100111;
            15'd17253: log10_cal = 16'b0000010011101000;
            15'd17254: log10_cal = 16'b0000010011101000;
            15'd17255: log10_cal = 16'b0000010011101000;
            15'd17256: log10_cal = 16'b0000010011101000;
            15'd17257: log10_cal = 16'b0000010011101000;
            15'd17258: log10_cal = 16'b0000010011101000;
            15'd17259: log10_cal = 16'b0000010011101000;
            15'd17260: log10_cal = 16'b0000010011101000;
            15'd17261: log10_cal = 16'b0000010011101000;
            15'd17262: log10_cal = 16'b0000010011101000;
            15'd17263: log10_cal = 16'b0000010011101000;
            15'd17264: log10_cal = 16'b0000010011101000;
            15'd17265: log10_cal = 16'b0000010011101000;
            15'd17266: log10_cal = 16'b0000010011101000;
            15'd17267: log10_cal = 16'b0000010011101000;
            15'd17268: log10_cal = 16'b0000010011101000;
            15'd17269: log10_cal = 16'b0000010011101000;
            15'd17270: log10_cal = 16'b0000010011101000;
            15'd17271: log10_cal = 16'b0000010011101000;
            15'd17272: log10_cal = 16'b0000010011101000;
            15'd17273: log10_cal = 16'b0000010011101000;
            15'd17274: log10_cal = 16'b0000010011101000;
            15'd17275: log10_cal = 16'b0000010011101000;
            15'd17276: log10_cal = 16'b0000010011101000;
            15'd17277: log10_cal = 16'b0000010011101000;
            15'd17278: log10_cal = 16'b0000010011101000;
            15'd17279: log10_cal = 16'b0000010011101000;
            15'd17280: log10_cal = 16'b0000010011101000;
            15'd17281: log10_cal = 16'b0000010011101000;
            15'd17282: log10_cal = 16'b0000010011101000;
            15'd17283: log10_cal = 16'b0000010011101000;
            15'd17284: log10_cal = 16'b0000010011101000;
            15'd17285: log10_cal = 16'b0000010011101000;
            15'd17286: log10_cal = 16'b0000010011101000;
            15'd17287: log10_cal = 16'b0000010011101000;
            15'd17288: log10_cal = 16'b0000010011101000;
            15'd17289: log10_cal = 16'b0000010011101000;
            15'd17290: log10_cal = 16'b0000010011101000;
            15'd17291: log10_cal = 16'b0000010011101000;
            15'd17292: log10_cal = 16'b0000010011101001;
            15'd17293: log10_cal = 16'b0000010011101001;
            15'd17294: log10_cal = 16'b0000010011101001;
            15'd17295: log10_cal = 16'b0000010011101001;
            15'd17296: log10_cal = 16'b0000010011101001;
            15'd17297: log10_cal = 16'b0000010011101001;
            15'd17298: log10_cal = 16'b0000010011101001;
            15'd17299: log10_cal = 16'b0000010011101001;
            15'd17300: log10_cal = 16'b0000010011101001;
            15'd17301: log10_cal = 16'b0000010011101001;
            15'd17302: log10_cal = 16'b0000010011101001;
            15'd17303: log10_cal = 16'b0000010011101001;
            15'd17304: log10_cal = 16'b0000010011101001;
            15'd17305: log10_cal = 16'b0000010011101001;
            15'd17306: log10_cal = 16'b0000010011101001;
            15'd17307: log10_cal = 16'b0000010011101001;
            15'd17308: log10_cal = 16'b0000010011101001;
            15'd17309: log10_cal = 16'b0000010011101001;
            15'd17310: log10_cal = 16'b0000010011101001;
            15'd17311: log10_cal = 16'b0000010011101001;
            15'd17312: log10_cal = 16'b0000010011101001;
            15'd17313: log10_cal = 16'b0000010011101001;
            15'd17314: log10_cal = 16'b0000010011101001;
            15'd17315: log10_cal = 16'b0000010011101001;
            15'd17316: log10_cal = 16'b0000010011101001;
            15'd17317: log10_cal = 16'b0000010011101001;
            15'd17318: log10_cal = 16'b0000010011101001;
            15'd17319: log10_cal = 16'b0000010011101001;
            15'd17320: log10_cal = 16'b0000010011101001;
            15'd17321: log10_cal = 16'b0000010011101001;
            15'd17322: log10_cal = 16'b0000010011101001;
            15'd17323: log10_cal = 16'b0000010011101001;
            15'd17324: log10_cal = 16'b0000010011101001;
            15'd17325: log10_cal = 16'b0000010011101001;
            15'd17326: log10_cal = 16'b0000010011101001;
            15'd17327: log10_cal = 16'b0000010011101001;
            15'd17328: log10_cal = 16'b0000010011101001;
            15'd17329: log10_cal = 16'b0000010011101001;
            15'd17330: log10_cal = 16'b0000010011101001;
            15'd17331: log10_cal = 16'b0000010011101010;
            15'd17332: log10_cal = 16'b0000010011101010;
            15'd17333: log10_cal = 16'b0000010011101010;
            15'd17334: log10_cal = 16'b0000010011101010;
            15'd17335: log10_cal = 16'b0000010011101010;
            15'd17336: log10_cal = 16'b0000010011101010;
            15'd17337: log10_cal = 16'b0000010011101010;
            15'd17338: log10_cal = 16'b0000010011101010;
            15'd17339: log10_cal = 16'b0000010011101010;
            15'd17340: log10_cal = 16'b0000010011101010;
            15'd17341: log10_cal = 16'b0000010011101010;
            15'd17342: log10_cal = 16'b0000010011101010;
            15'd17343: log10_cal = 16'b0000010011101010;
            15'd17344: log10_cal = 16'b0000010011101010;
            15'd17345: log10_cal = 16'b0000010011101010;
            15'd17346: log10_cal = 16'b0000010011101010;
            15'd17347: log10_cal = 16'b0000010011101010;
            15'd17348: log10_cal = 16'b0000010011101010;
            15'd17349: log10_cal = 16'b0000010011101010;
            15'd17350: log10_cal = 16'b0000010011101010;
            15'd17351: log10_cal = 16'b0000010011101010;
            15'd17352: log10_cal = 16'b0000010011101010;
            15'd17353: log10_cal = 16'b0000010011101010;
            15'd17354: log10_cal = 16'b0000010011101010;
            15'd17355: log10_cal = 16'b0000010011101010;
            15'd17356: log10_cal = 16'b0000010011101010;
            15'd17357: log10_cal = 16'b0000010011101010;
            15'd17358: log10_cal = 16'b0000010011101010;
            15'd17359: log10_cal = 16'b0000010011101010;
            15'd17360: log10_cal = 16'b0000010011101010;
            15'd17361: log10_cal = 16'b0000010011101010;
            15'd17362: log10_cal = 16'b0000010011101010;
            15'd17363: log10_cal = 16'b0000010011101010;
            15'd17364: log10_cal = 16'b0000010011101010;
            15'd17365: log10_cal = 16'b0000010011101010;
            15'd17366: log10_cal = 16'b0000010011101010;
            15'd17367: log10_cal = 16'b0000010011101010;
            15'd17368: log10_cal = 16'b0000010011101010;
            15'd17369: log10_cal = 16'b0000010011101010;
            15'd17370: log10_cal = 16'b0000010011101011;
            15'd17371: log10_cal = 16'b0000010011101011;
            15'd17372: log10_cal = 16'b0000010011101011;
            15'd17373: log10_cal = 16'b0000010011101011;
            15'd17374: log10_cal = 16'b0000010011101011;
            15'd17375: log10_cal = 16'b0000010011101011;
            15'd17376: log10_cal = 16'b0000010011101011;
            15'd17377: log10_cal = 16'b0000010011101011;
            15'd17378: log10_cal = 16'b0000010011101011;
            15'd17379: log10_cal = 16'b0000010011101011;
            15'd17380: log10_cal = 16'b0000010011101011;
            15'd17381: log10_cal = 16'b0000010011101011;
            15'd17382: log10_cal = 16'b0000010011101011;
            15'd17383: log10_cal = 16'b0000010011101011;
            15'd17384: log10_cal = 16'b0000010011101011;
            15'd17385: log10_cal = 16'b0000010011101011;
            15'd17386: log10_cal = 16'b0000010011101011;
            15'd17387: log10_cal = 16'b0000010011101011;
            15'd17388: log10_cal = 16'b0000010011101011;
            15'd17389: log10_cal = 16'b0000010011101011;
            15'd17390: log10_cal = 16'b0000010011101011;
            15'd17391: log10_cal = 16'b0000010011101011;
            15'd17392: log10_cal = 16'b0000010011101011;
            15'd17393: log10_cal = 16'b0000010011101011;
            15'd17394: log10_cal = 16'b0000010011101011;
            15'd17395: log10_cal = 16'b0000010011101011;
            15'd17396: log10_cal = 16'b0000010011101011;
            15'd17397: log10_cal = 16'b0000010011101011;
            15'd17398: log10_cal = 16'b0000010011101011;
            15'd17399: log10_cal = 16'b0000010011101011;
            15'd17400: log10_cal = 16'b0000010011101011;
            15'd17401: log10_cal = 16'b0000010011101011;
            15'd17402: log10_cal = 16'b0000010011101011;
            15'd17403: log10_cal = 16'b0000010011101011;
            15'd17404: log10_cal = 16'b0000010011101011;
            15'd17405: log10_cal = 16'b0000010011101011;
            15'd17406: log10_cal = 16'b0000010011101011;
            15'd17407: log10_cal = 16'b0000010011101011;
            15'd17408: log10_cal = 16'b0000010011101011;
            15'd17409: log10_cal = 16'b0000010011101100;
            15'd17410: log10_cal = 16'b0000010011101100;
            15'd17411: log10_cal = 16'b0000010011101100;
            15'd17412: log10_cal = 16'b0000010011101100;
            15'd17413: log10_cal = 16'b0000010011101100;
            15'd17414: log10_cal = 16'b0000010011101100;
            15'd17415: log10_cal = 16'b0000010011101100;
            15'd17416: log10_cal = 16'b0000010011101100;
            15'd17417: log10_cal = 16'b0000010011101100;
            15'd17418: log10_cal = 16'b0000010011101100;
            15'd17419: log10_cal = 16'b0000010011101100;
            15'd17420: log10_cal = 16'b0000010011101100;
            15'd17421: log10_cal = 16'b0000010011101100;
            15'd17422: log10_cal = 16'b0000010011101100;
            15'd17423: log10_cal = 16'b0000010011101100;
            15'd17424: log10_cal = 16'b0000010011101100;
            15'd17425: log10_cal = 16'b0000010011101100;
            15'd17426: log10_cal = 16'b0000010011101100;
            15'd17427: log10_cal = 16'b0000010011101100;
            15'd17428: log10_cal = 16'b0000010011101100;
            15'd17429: log10_cal = 16'b0000010011101100;
            15'd17430: log10_cal = 16'b0000010011101100;
            15'd17431: log10_cal = 16'b0000010011101100;
            15'd17432: log10_cal = 16'b0000010011101100;
            15'd17433: log10_cal = 16'b0000010011101100;
            15'd17434: log10_cal = 16'b0000010011101100;
            15'd17435: log10_cal = 16'b0000010011101100;
            15'd17436: log10_cal = 16'b0000010011101100;
            15'd17437: log10_cal = 16'b0000010011101100;
            15'd17438: log10_cal = 16'b0000010011101100;
            15'd17439: log10_cal = 16'b0000010011101100;
            15'd17440: log10_cal = 16'b0000010011101100;
            15'd17441: log10_cal = 16'b0000010011101100;
            15'd17442: log10_cal = 16'b0000010011101100;
            15'd17443: log10_cal = 16'b0000010011101100;
            15'd17444: log10_cal = 16'b0000010011101100;
            15'd17445: log10_cal = 16'b0000010011101100;
            15'd17446: log10_cal = 16'b0000010011101100;
            15'd17447: log10_cal = 16'b0000010011101100;
            15'd17448: log10_cal = 16'b0000010011101101;
            15'd17449: log10_cal = 16'b0000010011101101;
            15'd17450: log10_cal = 16'b0000010011101101;
            15'd17451: log10_cal = 16'b0000010011101101;
            15'd17452: log10_cal = 16'b0000010011101101;
            15'd17453: log10_cal = 16'b0000010011101101;
            15'd17454: log10_cal = 16'b0000010011101101;
            15'd17455: log10_cal = 16'b0000010011101101;
            15'd17456: log10_cal = 16'b0000010011101101;
            15'd17457: log10_cal = 16'b0000010011101101;
            15'd17458: log10_cal = 16'b0000010011101101;
            15'd17459: log10_cal = 16'b0000010011101101;
            15'd17460: log10_cal = 16'b0000010011101101;
            15'd17461: log10_cal = 16'b0000010011101101;
            15'd17462: log10_cal = 16'b0000010011101101;
            15'd17463: log10_cal = 16'b0000010011101101;
            15'd17464: log10_cal = 16'b0000010011101101;
            15'd17465: log10_cal = 16'b0000010011101101;
            15'd17466: log10_cal = 16'b0000010011101101;
            15'd17467: log10_cal = 16'b0000010011101101;
            15'd17468: log10_cal = 16'b0000010011101101;
            15'd17469: log10_cal = 16'b0000010011101101;
            15'd17470: log10_cal = 16'b0000010011101101;
            15'd17471: log10_cal = 16'b0000010011101101;
            15'd17472: log10_cal = 16'b0000010011101101;
            15'd17473: log10_cal = 16'b0000010011101101;
            15'd17474: log10_cal = 16'b0000010011101101;
            15'd17475: log10_cal = 16'b0000010011101101;
            15'd17476: log10_cal = 16'b0000010011101101;
            15'd17477: log10_cal = 16'b0000010011101101;
            15'd17478: log10_cal = 16'b0000010011101101;
            15'd17479: log10_cal = 16'b0000010011101101;
            15'd17480: log10_cal = 16'b0000010011101101;
            15'd17481: log10_cal = 16'b0000010011101101;
            15'd17482: log10_cal = 16'b0000010011101101;
            15'd17483: log10_cal = 16'b0000010011101101;
            15'd17484: log10_cal = 16'b0000010011101101;
            15'd17485: log10_cal = 16'b0000010011101101;
            15'd17486: log10_cal = 16'b0000010011101101;
            15'd17487: log10_cal = 16'b0000010011101101;
            15'd17488: log10_cal = 16'b0000010011101110;
            15'd17489: log10_cal = 16'b0000010011101110;
            15'd17490: log10_cal = 16'b0000010011101110;
            15'd17491: log10_cal = 16'b0000010011101110;
            15'd17492: log10_cal = 16'b0000010011101110;
            15'd17493: log10_cal = 16'b0000010011101110;
            15'd17494: log10_cal = 16'b0000010011101110;
            15'd17495: log10_cal = 16'b0000010011101110;
            15'd17496: log10_cal = 16'b0000010011101110;
            15'd17497: log10_cal = 16'b0000010011101110;
            15'd17498: log10_cal = 16'b0000010011101110;
            15'd17499: log10_cal = 16'b0000010011101110;
            15'd17500: log10_cal = 16'b0000010011101110;
            15'd17501: log10_cal = 16'b0000010011101110;
            15'd17502: log10_cal = 16'b0000010011101110;
            15'd17503: log10_cal = 16'b0000010011101110;
            15'd17504: log10_cal = 16'b0000010011101110;
            15'd17505: log10_cal = 16'b0000010011101110;
            15'd17506: log10_cal = 16'b0000010011101110;
            15'd17507: log10_cal = 16'b0000010011101110;
            15'd17508: log10_cal = 16'b0000010011101110;
            15'd17509: log10_cal = 16'b0000010011101110;
            15'd17510: log10_cal = 16'b0000010011101110;
            15'd17511: log10_cal = 16'b0000010011101110;
            15'd17512: log10_cal = 16'b0000010011101110;
            15'd17513: log10_cal = 16'b0000010011101110;
            15'd17514: log10_cal = 16'b0000010011101110;
            15'd17515: log10_cal = 16'b0000010011101110;
            15'd17516: log10_cal = 16'b0000010011101110;
            15'd17517: log10_cal = 16'b0000010011101110;
            15'd17518: log10_cal = 16'b0000010011101110;
            15'd17519: log10_cal = 16'b0000010011101110;
            15'd17520: log10_cal = 16'b0000010011101110;
            15'd17521: log10_cal = 16'b0000010011101110;
            15'd17522: log10_cal = 16'b0000010011101110;
            15'd17523: log10_cal = 16'b0000010011101110;
            15'd17524: log10_cal = 16'b0000010011101110;
            15'd17525: log10_cal = 16'b0000010011101110;
            15'd17526: log10_cal = 16'b0000010011101110;
            15'd17527: log10_cal = 16'b0000010011101111;
            15'd17528: log10_cal = 16'b0000010011101111;
            15'd17529: log10_cal = 16'b0000010011101111;
            15'd17530: log10_cal = 16'b0000010011101111;
            15'd17531: log10_cal = 16'b0000010011101111;
            15'd17532: log10_cal = 16'b0000010011101111;
            15'd17533: log10_cal = 16'b0000010011101111;
            15'd17534: log10_cal = 16'b0000010011101111;
            15'd17535: log10_cal = 16'b0000010011101111;
            15'd17536: log10_cal = 16'b0000010011101111;
            15'd17537: log10_cal = 16'b0000010011101111;
            15'd17538: log10_cal = 16'b0000010011101111;
            15'd17539: log10_cal = 16'b0000010011101111;
            15'd17540: log10_cal = 16'b0000010011101111;
            15'd17541: log10_cal = 16'b0000010011101111;
            15'd17542: log10_cal = 16'b0000010011101111;
            15'd17543: log10_cal = 16'b0000010011101111;
            15'd17544: log10_cal = 16'b0000010011101111;
            15'd17545: log10_cal = 16'b0000010011101111;
            15'd17546: log10_cal = 16'b0000010011101111;
            15'd17547: log10_cal = 16'b0000010011101111;
            15'd17548: log10_cal = 16'b0000010011101111;
            15'd17549: log10_cal = 16'b0000010011101111;
            15'd17550: log10_cal = 16'b0000010011101111;
            15'd17551: log10_cal = 16'b0000010011101111;
            15'd17552: log10_cal = 16'b0000010011101111;
            15'd17553: log10_cal = 16'b0000010011101111;
            15'd17554: log10_cal = 16'b0000010011101111;
            15'd17555: log10_cal = 16'b0000010011101111;
            15'd17556: log10_cal = 16'b0000010011101111;
            15'd17557: log10_cal = 16'b0000010011101111;
            15'd17558: log10_cal = 16'b0000010011101111;
            15'd17559: log10_cal = 16'b0000010011101111;
            15'd17560: log10_cal = 16'b0000010011101111;
            15'd17561: log10_cal = 16'b0000010011101111;
            15'd17562: log10_cal = 16'b0000010011101111;
            15'd17563: log10_cal = 16'b0000010011101111;
            15'd17564: log10_cal = 16'b0000010011101111;
            15'd17565: log10_cal = 16'b0000010011101111;
            15'd17566: log10_cal = 16'b0000010011101111;
            15'd17567: log10_cal = 16'b0000010011110000;
            15'd17568: log10_cal = 16'b0000010011110000;
            15'd17569: log10_cal = 16'b0000010011110000;
            15'd17570: log10_cal = 16'b0000010011110000;
            15'd17571: log10_cal = 16'b0000010011110000;
            15'd17572: log10_cal = 16'b0000010011110000;
            15'd17573: log10_cal = 16'b0000010011110000;
            15'd17574: log10_cal = 16'b0000010011110000;
            15'd17575: log10_cal = 16'b0000010011110000;
            15'd17576: log10_cal = 16'b0000010011110000;
            15'd17577: log10_cal = 16'b0000010011110000;
            15'd17578: log10_cal = 16'b0000010011110000;
            15'd17579: log10_cal = 16'b0000010011110000;
            15'd17580: log10_cal = 16'b0000010011110000;
            15'd17581: log10_cal = 16'b0000010011110000;
            15'd17582: log10_cal = 16'b0000010011110000;
            15'd17583: log10_cal = 16'b0000010011110000;
            15'd17584: log10_cal = 16'b0000010011110000;
            15'd17585: log10_cal = 16'b0000010011110000;
            15'd17586: log10_cal = 16'b0000010011110000;
            15'd17587: log10_cal = 16'b0000010011110000;
            15'd17588: log10_cal = 16'b0000010011110000;
            15'd17589: log10_cal = 16'b0000010011110000;
            15'd17590: log10_cal = 16'b0000010011110000;
            15'd17591: log10_cal = 16'b0000010011110000;
            15'd17592: log10_cal = 16'b0000010011110000;
            15'd17593: log10_cal = 16'b0000010011110000;
            15'd17594: log10_cal = 16'b0000010011110000;
            15'd17595: log10_cal = 16'b0000010011110000;
            15'd17596: log10_cal = 16'b0000010011110000;
            15'd17597: log10_cal = 16'b0000010011110000;
            15'd17598: log10_cal = 16'b0000010011110000;
            15'd17599: log10_cal = 16'b0000010011110000;
            15'd17600: log10_cal = 16'b0000010011110000;
            15'd17601: log10_cal = 16'b0000010011110000;
            15'd17602: log10_cal = 16'b0000010011110000;
            15'd17603: log10_cal = 16'b0000010011110000;
            15'd17604: log10_cal = 16'b0000010011110000;
            15'd17605: log10_cal = 16'b0000010011110000;
            15'd17606: log10_cal = 16'b0000010011110001;
            15'd17607: log10_cal = 16'b0000010011110001;
            15'd17608: log10_cal = 16'b0000010011110001;
            15'd17609: log10_cal = 16'b0000010011110001;
            15'd17610: log10_cal = 16'b0000010011110001;
            15'd17611: log10_cal = 16'b0000010011110001;
            15'd17612: log10_cal = 16'b0000010011110001;
            15'd17613: log10_cal = 16'b0000010011110001;
            15'd17614: log10_cal = 16'b0000010011110001;
            15'd17615: log10_cal = 16'b0000010011110001;
            15'd17616: log10_cal = 16'b0000010011110001;
            15'd17617: log10_cal = 16'b0000010011110001;
            15'd17618: log10_cal = 16'b0000010011110001;
            15'd17619: log10_cal = 16'b0000010011110001;
            15'd17620: log10_cal = 16'b0000010011110001;
            15'd17621: log10_cal = 16'b0000010011110001;
            15'd17622: log10_cal = 16'b0000010011110001;
            15'd17623: log10_cal = 16'b0000010011110001;
            15'd17624: log10_cal = 16'b0000010011110001;
            15'd17625: log10_cal = 16'b0000010011110001;
            15'd17626: log10_cal = 16'b0000010011110001;
            15'd17627: log10_cal = 16'b0000010011110001;
            15'd17628: log10_cal = 16'b0000010011110001;
            15'd17629: log10_cal = 16'b0000010011110001;
            15'd17630: log10_cal = 16'b0000010011110001;
            15'd17631: log10_cal = 16'b0000010011110001;
            15'd17632: log10_cal = 16'b0000010011110001;
            15'd17633: log10_cal = 16'b0000010011110001;
            15'd17634: log10_cal = 16'b0000010011110001;
            15'd17635: log10_cal = 16'b0000010011110001;
            15'd17636: log10_cal = 16'b0000010011110001;
            15'd17637: log10_cal = 16'b0000010011110001;
            15'd17638: log10_cal = 16'b0000010011110001;
            15'd17639: log10_cal = 16'b0000010011110001;
            15'd17640: log10_cal = 16'b0000010011110001;
            15'd17641: log10_cal = 16'b0000010011110001;
            15'd17642: log10_cal = 16'b0000010011110001;
            15'd17643: log10_cal = 16'b0000010011110001;
            15'd17644: log10_cal = 16'b0000010011110001;
            15'd17645: log10_cal = 16'b0000010011110001;
            15'd17646: log10_cal = 16'b0000010011110010;
            15'd17647: log10_cal = 16'b0000010011110010;
            15'd17648: log10_cal = 16'b0000010011110010;
            15'd17649: log10_cal = 16'b0000010011110010;
            15'd17650: log10_cal = 16'b0000010011110010;
            15'd17651: log10_cal = 16'b0000010011110010;
            15'd17652: log10_cal = 16'b0000010011110010;
            15'd17653: log10_cal = 16'b0000010011110010;
            15'd17654: log10_cal = 16'b0000010011110010;
            15'd17655: log10_cal = 16'b0000010011110010;
            15'd17656: log10_cal = 16'b0000010011110010;
            15'd17657: log10_cal = 16'b0000010011110010;
            15'd17658: log10_cal = 16'b0000010011110010;
            15'd17659: log10_cal = 16'b0000010011110010;
            15'd17660: log10_cal = 16'b0000010011110010;
            15'd17661: log10_cal = 16'b0000010011110010;
            15'd17662: log10_cal = 16'b0000010011110010;
            15'd17663: log10_cal = 16'b0000010011110010;
            15'd17664: log10_cal = 16'b0000010011110010;
            15'd17665: log10_cal = 16'b0000010011110010;
            15'd17666: log10_cal = 16'b0000010011110010;
            15'd17667: log10_cal = 16'b0000010011110010;
            15'd17668: log10_cal = 16'b0000010011110010;
            15'd17669: log10_cal = 16'b0000010011110010;
            15'd17670: log10_cal = 16'b0000010011110010;
            15'd17671: log10_cal = 16'b0000010011110010;
            15'd17672: log10_cal = 16'b0000010011110010;
            15'd17673: log10_cal = 16'b0000010011110010;
            15'd17674: log10_cal = 16'b0000010011110010;
            15'd17675: log10_cal = 16'b0000010011110010;
            15'd17676: log10_cal = 16'b0000010011110010;
            15'd17677: log10_cal = 16'b0000010011110010;
            15'd17678: log10_cal = 16'b0000010011110010;
            15'd17679: log10_cal = 16'b0000010011110010;
            15'd17680: log10_cal = 16'b0000010011110010;
            15'd17681: log10_cal = 16'b0000010011110010;
            15'd17682: log10_cal = 16'b0000010011110010;
            15'd17683: log10_cal = 16'b0000010011110010;
            15'd17684: log10_cal = 16'b0000010011110010;
            15'd17685: log10_cal = 16'b0000010011110011;
            15'd17686: log10_cal = 16'b0000010011110011;
            15'd17687: log10_cal = 16'b0000010011110011;
            15'd17688: log10_cal = 16'b0000010011110011;
            15'd17689: log10_cal = 16'b0000010011110011;
            15'd17690: log10_cal = 16'b0000010011110011;
            15'd17691: log10_cal = 16'b0000010011110011;
            15'd17692: log10_cal = 16'b0000010011110011;
            15'd17693: log10_cal = 16'b0000010011110011;
            15'd17694: log10_cal = 16'b0000010011110011;
            15'd17695: log10_cal = 16'b0000010011110011;
            15'd17696: log10_cal = 16'b0000010011110011;
            15'd17697: log10_cal = 16'b0000010011110011;
            15'd17698: log10_cal = 16'b0000010011110011;
            15'd17699: log10_cal = 16'b0000010011110011;
            15'd17700: log10_cal = 16'b0000010011110011;
            15'd17701: log10_cal = 16'b0000010011110011;
            15'd17702: log10_cal = 16'b0000010011110011;
            15'd17703: log10_cal = 16'b0000010011110011;
            15'd17704: log10_cal = 16'b0000010011110011;
            15'd17705: log10_cal = 16'b0000010011110011;
            15'd17706: log10_cal = 16'b0000010011110011;
            15'd17707: log10_cal = 16'b0000010011110011;
            15'd17708: log10_cal = 16'b0000010011110011;
            15'd17709: log10_cal = 16'b0000010011110011;
            15'd17710: log10_cal = 16'b0000010011110011;
            15'd17711: log10_cal = 16'b0000010011110011;
            15'd17712: log10_cal = 16'b0000010011110011;
            15'd17713: log10_cal = 16'b0000010011110011;
            15'd17714: log10_cal = 16'b0000010011110011;
            15'd17715: log10_cal = 16'b0000010011110011;
            15'd17716: log10_cal = 16'b0000010011110011;
            15'd17717: log10_cal = 16'b0000010011110011;
            15'd17718: log10_cal = 16'b0000010011110011;
            15'd17719: log10_cal = 16'b0000010011110011;
            15'd17720: log10_cal = 16'b0000010011110011;
            15'd17721: log10_cal = 16'b0000010011110011;
            15'd17722: log10_cal = 16'b0000010011110011;
            15'd17723: log10_cal = 16'b0000010011110011;
            15'd17724: log10_cal = 16'b0000010011110011;
            15'd17725: log10_cal = 16'b0000010011110100;
            15'd17726: log10_cal = 16'b0000010011110100;
            15'd17727: log10_cal = 16'b0000010011110100;
            15'd17728: log10_cal = 16'b0000010011110100;
            15'd17729: log10_cal = 16'b0000010011110100;
            15'd17730: log10_cal = 16'b0000010011110100;
            15'd17731: log10_cal = 16'b0000010011110100;
            15'd17732: log10_cal = 16'b0000010011110100;
            15'd17733: log10_cal = 16'b0000010011110100;
            15'd17734: log10_cal = 16'b0000010011110100;
            15'd17735: log10_cal = 16'b0000010011110100;
            15'd17736: log10_cal = 16'b0000010011110100;
            15'd17737: log10_cal = 16'b0000010011110100;
            15'd17738: log10_cal = 16'b0000010011110100;
            15'd17739: log10_cal = 16'b0000010011110100;
            15'd17740: log10_cal = 16'b0000010011110100;
            15'd17741: log10_cal = 16'b0000010011110100;
            15'd17742: log10_cal = 16'b0000010011110100;
            15'd17743: log10_cal = 16'b0000010011110100;
            15'd17744: log10_cal = 16'b0000010011110100;
            15'd17745: log10_cal = 16'b0000010011110100;
            15'd17746: log10_cal = 16'b0000010011110100;
            15'd17747: log10_cal = 16'b0000010011110100;
            15'd17748: log10_cal = 16'b0000010011110100;
            15'd17749: log10_cal = 16'b0000010011110100;
            15'd17750: log10_cal = 16'b0000010011110100;
            15'd17751: log10_cal = 16'b0000010011110100;
            15'd17752: log10_cal = 16'b0000010011110100;
            15'd17753: log10_cal = 16'b0000010011110100;
            15'd17754: log10_cal = 16'b0000010011110100;
            15'd17755: log10_cal = 16'b0000010011110100;
            15'd17756: log10_cal = 16'b0000010011110100;
            15'd17757: log10_cal = 16'b0000010011110100;
            15'd17758: log10_cal = 16'b0000010011110100;
            15'd17759: log10_cal = 16'b0000010011110100;
            15'd17760: log10_cal = 16'b0000010011110100;
            15'd17761: log10_cal = 16'b0000010011110100;
            15'd17762: log10_cal = 16'b0000010011110100;
            15'd17763: log10_cal = 16'b0000010011110100;
            15'd17764: log10_cal = 16'b0000010011110100;
            15'd17765: log10_cal = 16'b0000010011110101;
            15'd17766: log10_cal = 16'b0000010011110101;
            15'd17767: log10_cal = 16'b0000010011110101;
            15'd17768: log10_cal = 16'b0000010011110101;
            15'd17769: log10_cal = 16'b0000010011110101;
            15'd17770: log10_cal = 16'b0000010011110101;
            15'd17771: log10_cal = 16'b0000010011110101;
            15'd17772: log10_cal = 16'b0000010011110101;
            15'd17773: log10_cal = 16'b0000010011110101;
            15'd17774: log10_cal = 16'b0000010011110101;
            15'd17775: log10_cal = 16'b0000010011110101;
            15'd17776: log10_cal = 16'b0000010011110101;
            15'd17777: log10_cal = 16'b0000010011110101;
            15'd17778: log10_cal = 16'b0000010011110101;
            15'd17779: log10_cal = 16'b0000010011110101;
            15'd17780: log10_cal = 16'b0000010011110101;
            15'd17781: log10_cal = 16'b0000010011110101;
            15'd17782: log10_cal = 16'b0000010011110101;
            15'd17783: log10_cal = 16'b0000010011110101;
            15'd17784: log10_cal = 16'b0000010011110101;
            15'd17785: log10_cal = 16'b0000010011110101;
            15'd17786: log10_cal = 16'b0000010011110101;
            15'd17787: log10_cal = 16'b0000010011110101;
            15'd17788: log10_cal = 16'b0000010011110101;
            15'd17789: log10_cal = 16'b0000010011110101;
            15'd17790: log10_cal = 16'b0000010011110101;
            15'd17791: log10_cal = 16'b0000010011110101;
            15'd17792: log10_cal = 16'b0000010011110101;
            15'd17793: log10_cal = 16'b0000010011110101;
            15'd17794: log10_cal = 16'b0000010011110101;
            15'd17795: log10_cal = 16'b0000010011110101;
            15'd17796: log10_cal = 16'b0000010011110101;
            15'd17797: log10_cal = 16'b0000010011110101;
            15'd17798: log10_cal = 16'b0000010011110101;
            15'd17799: log10_cal = 16'b0000010011110101;
            15'd17800: log10_cal = 16'b0000010011110101;
            15'd17801: log10_cal = 16'b0000010011110101;
            15'd17802: log10_cal = 16'b0000010011110101;
            15'd17803: log10_cal = 16'b0000010011110101;
            15'd17804: log10_cal = 16'b0000010011110101;
            15'd17805: log10_cal = 16'b0000010011110110;
            15'd17806: log10_cal = 16'b0000010011110110;
            15'd17807: log10_cal = 16'b0000010011110110;
            15'd17808: log10_cal = 16'b0000010011110110;
            15'd17809: log10_cal = 16'b0000010011110110;
            15'd17810: log10_cal = 16'b0000010011110110;
            15'd17811: log10_cal = 16'b0000010011110110;
            15'd17812: log10_cal = 16'b0000010011110110;
            15'd17813: log10_cal = 16'b0000010011110110;
            15'd17814: log10_cal = 16'b0000010011110110;
            15'd17815: log10_cal = 16'b0000010011110110;
            15'd17816: log10_cal = 16'b0000010011110110;
            15'd17817: log10_cal = 16'b0000010011110110;
            15'd17818: log10_cal = 16'b0000010011110110;
            15'd17819: log10_cal = 16'b0000010011110110;
            15'd17820: log10_cal = 16'b0000010011110110;
            15'd17821: log10_cal = 16'b0000010011110110;
            15'd17822: log10_cal = 16'b0000010011110110;
            15'd17823: log10_cal = 16'b0000010011110110;
            15'd17824: log10_cal = 16'b0000010011110110;
            15'd17825: log10_cal = 16'b0000010011110110;
            15'd17826: log10_cal = 16'b0000010011110110;
            15'd17827: log10_cal = 16'b0000010011110110;
            15'd17828: log10_cal = 16'b0000010011110110;
            15'd17829: log10_cal = 16'b0000010011110110;
            15'd17830: log10_cal = 16'b0000010011110110;
            15'd17831: log10_cal = 16'b0000010011110110;
            15'd17832: log10_cal = 16'b0000010011110110;
            15'd17833: log10_cal = 16'b0000010011110110;
            15'd17834: log10_cal = 16'b0000010011110110;
            15'd17835: log10_cal = 16'b0000010011110110;
            15'd17836: log10_cal = 16'b0000010011110110;
            15'd17837: log10_cal = 16'b0000010011110110;
            15'd17838: log10_cal = 16'b0000010011110110;
            15'd17839: log10_cal = 16'b0000010011110110;
            15'd17840: log10_cal = 16'b0000010011110110;
            15'd17841: log10_cal = 16'b0000010011110110;
            15'd17842: log10_cal = 16'b0000010011110110;
            15'd17843: log10_cal = 16'b0000010011110110;
            15'd17844: log10_cal = 16'b0000010011110110;
            15'd17845: log10_cal = 16'b0000010011110111;
            15'd17846: log10_cal = 16'b0000010011110111;
            15'd17847: log10_cal = 16'b0000010011110111;
            15'd17848: log10_cal = 16'b0000010011110111;
            15'd17849: log10_cal = 16'b0000010011110111;
            15'd17850: log10_cal = 16'b0000010011110111;
            15'd17851: log10_cal = 16'b0000010011110111;
            15'd17852: log10_cal = 16'b0000010011110111;
            15'd17853: log10_cal = 16'b0000010011110111;
            15'd17854: log10_cal = 16'b0000010011110111;
            15'd17855: log10_cal = 16'b0000010011110111;
            15'd17856: log10_cal = 16'b0000010011110111;
            15'd17857: log10_cal = 16'b0000010011110111;
            15'd17858: log10_cal = 16'b0000010011110111;
            15'd17859: log10_cal = 16'b0000010011110111;
            15'd17860: log10_cal = 16'b0000010011110111;
            15'd17861: log10_cal = 16'b0000010011110111;
            15'd17862: log10_cal = 16'b0000010011110111;
            15'd17863: log10_cal = 16'b0000010011110111;
            15'd17864: log10_cal = 16'b0000010011110111;
            15'd17865: log10_cal = 16'b0000010011110111;
            15'd17866: log10_cal = 16'b0000010011110111;
            15'd17867: log10_cal = 16'b0000010011110111;
            15'd17868: log10_cal = 16'b0000010011110111;
            15'd17869: log10_cal = 16'b0000010011110111;
            15'd17870: log10_cal = 16'b0000010011110111;
            15'd17871: log10_cal = 16'b0000010011110111;
            15'd17872: log10_cal = 16'b0000010011110111;
            15'd17873: log10_cal = 16'b0000010011110111;
            15'd17874: log10_cal = 16'b0000010011110111;
            15'd17875: log10_cal = 16'b0000010011110111;
            15'd17876: log10_cal = 16'b0000010011110111;
            15'd17877: log10_cal = 16'b0000010011110111;
            15'd17878: log10_cal = 16'b0000010011110111;
            15'd17879: log10_cal = 16'b0000010011110111;
            15'd17880: log10_cal = 16'b0000010011110111;
            15'd17881: log10_cal = 16'b0000010011110111;
            15'd17882: log10_cal = 16'b0000010011110111;
            15'd17883: log10_cal = 16'b0000010011110111;
            15'd17884: log10_cal = 16'b0000010011110111;
            15'd17885: log10_cal = 16'b0000010011111000;
            15'd17886: log10_cal = 16'b0000010011111000;
            15'd17887: log10_cal = 16'b0000010011111000;
            15'd17888: log10_cal = 16'b0000010011111000;
            15'd17889: log10_cal = 16'b0000010011111000;
            15'd17890: log10_cal = 16'b0000010011111000;
            15'd17891: log10_cal = 16'b0000010011111000;
            15'd17892: log10_cal = 16'b0000010011111000;
            15'd17893: log10_cal = 16'b0000010011111000;
            15'd17894: log10_cal = 16'b0000010011111000;
            15'd17895: log10_cal = 16'b0000010011111000;
            15'd17896: log10_cal = 16'b0000010011111000;
            15'd17897: log10_cal = 16'b0000010011111000;
            15'd17898: log10_cal = 16'b0000010011111000;
            15'd17899: log10_cal = 16'b0000010011111000;
            15'd17900: log10_cal = 16'b0000010011111000;
            15'd17901: log10_cal = 16'b0000010011111000;
            15'd17902: log10_cal = 16'b0000010011111000;
            15'd17903: log10_cal = 16'b0000010011111000;
            15'd17904: log10_cal = 16'b0000010011111000;
            15'd17905: log10_cal = 16'b0000010011111000;
            15'd17906: log10_cal = 16'b0000010011111000;
            15'd17907: log10_cal = 16'b0000010011111000;
            15'd17908: log10_cal = 16'b0000010011111000;
            15'd17909: log10_cal = 16'b0000010011111000;
            15'd17910: log10_cal = 16'b0000010011111000;
            15'd17911: log10_cal = 16'b0000010011111000;
            15'd17912: log10_cal = 16'b0000010011111000;
            15'd17913: log10_cal = 16'b0000010011111000;
            15'd17914: log10_cal = 16'b0000010011111000;
            15'd17915: log10_cal = 16'b0000010011111000;
            15'd17916: log10_cal = 16'b0000010011111000;
            15'd17917: log10_cal = 16'b0000010011111000;
            15'd17918: log10_cal = 16'b0000010011111000;
            15'd17919: log10_cal = 16'b0000010011111000;
            15'd17920: log10_cal = 16'b0000010011111000;
            15'd17921: log10_cal = 16'b0000010011111000;
            15'd17922: log10_cal = 16'b0000010011111000;
            15'd17923: log10_cal = 16'b0000010011111000;
            15'd17924: log10_cal = 16'b0000010011111000;
            15'd17925: log10_cal = 16'b0000010011111000;
            15'd17926: log10_cal = 16'b0000010011111001;
            15'd17927: log10_cal = 16'b0000010011111001;
            15'd17928: log10_cal = 16'b0000010011111001;
            15'd17929: log10_cal = 16'b0000010011111001;
            15'd17930: log10_cal = 16'b0000010011111001;
            15'd17931: log10_cal = 16'b0000010011111001;
            15'd17932: log10_cal = 16'b0000010011111001;
            15'd17933: log10_cal = 16'b0000010011111001;
            15'd17934: log10_cal = 16'b0000010011111001;
            15'd17935: log10_cal = 16'b0000010011111001;
            15'd17936: log10_cal = 16'b0000010011111001;
            15'd17937: log10_cal = 16'b0000010011111001;
            15'd17938: log10_cal = 16'b0000010011111001;
            15'd17939: log10_cal = 16'b0000010011111001;
            15'd17940: log10_cal = 16'b0000010011111001;
            15'd17941: log10_cal = 16'b0000010011111001;
            15'd17942: log10_cal = 16'b0000010011111001;
            15'd17943: log10_cal = 16'b0000010011111001;
            15'd17944: log10_cal = 16'b0000010011111001;
            15'd17945: log10_cal = 16'b0000010011111001;
            15'd17946: log10_cal = 16'b0000010011111001;
            15'd17947: log10_cal = 16'b0000010011111001;
            15'd17948: log10_cal = 16'b0000010011111001;
            15'd17949: log10_cal = 16'b0000010011111001;
            15'd17950: log10_cal = 16'b0000010011111001;
            15'd17951: log10_cal = 16'b0000010011111001;
            15'd17952: log10_cal = 16'b0000010011111001;
            15'd17953: log10_cal = 16'b0000010011111001;
            15'd17954: log10_cal = 16'b0000010011111001;
            15'd17955: log10_cal = 16'b0000010011111001;
            15'd17956: log10_cal = 16'b0000010011111001;
            15'd17957: log10_cal = 16'b0000010011111001;
            15'd17958: log10_cal = 16'b0000010011111001;
            15'd17959: log10_cal = 16'b0000010011111001;
            15'd17960: log10_cal = 16'b0000010011111001;
            15'd17961: log10_cal = 16'b0000010011111001;
            15'd17962: log10_cal = 16'b0000010011111001;
            15'd17963: log10_cal = 16'b0000010011111001;
            15'd17964: log10_cal = 16'b0000010011111001;
            15'd17965: log10_cal = 16'b0000010011111001;
            15'd17966: log10_cal = 16'b0000010011111010;
            15'd17967: log10_cal = 16'b0000010011111010;
            15'd17968: log10_cal = 16'b0000010011111010;
            15'd17969: log10_cal = 16'b0000010011111010;
            15'd17970: log10_cal = 16'b0000010011111010;
            15'd17971: log10_cal = 16'b0000010011111010;
            15'd17972: log10_cal = 16'b0000010011111010;
            15'd17973: log10_cal = 16'b0000010011111010;
            15'd17974: log10_cal = 16'b0000010011111010;
            15'd17975: log10_cal = 16'b0000010011111010;
            15'd17976: log10_cal = 16'b0000010011111010;
            15'd17977: log10_cal = 16'b0000010011111010;
            15'd17978: log10_cal = 16'b0000010011111010;
            15'd17979: log10_cal = 16'b0000010011111010;
            15'd17980: log10_cal = 16'b0000010011111010;
            15'd17981: log10_cal = 16'b0000010011111010;
            15'd17982: log10_cal = 16'b0000010011111010;
            15'd17983: log10_cal = 16'b0000010011111010;
            15'd17984: log10_cal = 16'b0000010011111010;
            15'd17985: log10_cal = 16'b0000010011111010;
            15'd17986: log10_cal = 16'b0000010011111010;
            15'd17987: log10_cal = 16'b0000010011111010;
            15'd17988: log10_cal = 16'b0000010011111010;
            15'd17989: log10_cal = 16'b0000010011111010;
            15'd17990: log10_cal = 16'b0000010011111010;
            15'd17991: log10_cal = 16'b0000010011111010;
            15'd17992: log10_cal = 16'b0000010011111010;
            15'd17993: log10_cal = 16'b0000010011111010;
            15'd17994: log10_cal = 16'b0000010011111010;
            15'd17995: log10_cal = 16'b0000010011111010;
            15'd17996: log10_cal = 16'b0000010011111010;
            15'd17997: log10_cal = 16'b0000010011111010;
            15'd17998: log10_cal = 16'b0000010011111010;
            15'd17999: log10_cal = 16'b0000010011111010;
            15'd18000: log10_cal = 16'b0000010011111010;
            15'd18001: log10_cal = 16'b0000010011111010;
            15'd18002: log10_cal = 16'b0000010011111010;
            15'd18003: log10_cal = 16'b0000010011111010;
            15'd18004: log10_cal = 16'b0000010011111010;
            15'd18005: log10_cal = 16'b0000010011111010;
            15'd18006: log10_cal = 16'b0000010011111011;
            15'd18007: log10_cal = 16'b0000010011111011;
            15'd18008: log10_cal = 16'b0000010011111011;
            15'd18009: log10_cal = 16'b0000010011111011;
            15'd18010: log10_cal = 16'b0000010011111011;
            15'd18011: log10_cal = 16'b0000010011111011;
            15'd18012: log10_cal = 16'b0000010011111011;
            15'd18013: log10_cal = 16'b0000010011111011;
            15'd18014: log10_cal = 16'b0000010011111011;
            15'd18015: log10_cal = 16'b0000010011111011;
            15'd18016: log10_cal = 16'b0000010011111011;
            15'd18017: log10_cal = 16'b0000010011111011;
            15'd18018: log10_cal = 16'b0000010011111011;
            15'd18019: log10_cal = 16'b0000010011111011;
            15'd18020: log10_cal = 16'b0000010011111011;
            15'd18021: log10_cal = 16'b0000010011111011;
            15'd18022: log10_cal = 16'b0000010011111011;
            15'd18023: log10_cal = 16'b0000010011111011;
            15'd18024: log10_cal = 16'b0000010011111011;
            15'd18025: log10_cal = 16'b0000010011111011;
            15'd18026: log10_cal = 16'b0000010011111011;
            15'd18027: log10_cal = 16'b0000010011111011;
            15'd18028: log10_cal = 16'b0000010011111011;
            15'd18029: log10_cal = 16'b0000010011111011;
            15'd18030: log10_cal = 16'b0000010011111011;
            15'd18031: log10_cal = 16'b0000010011111011;
            15'd18032: log10_cal = 16'b0000010011111011;
            15'd18033: log10_cal = 16'b0000010011111011;
            15'd18034: log10_cal = 16'b0000010011111011;
            15'd18035: log10_cal = 16'b0000010011111011;
            15'd18036: log10_cal = 16'b0000010011111011;
            15'd18037: log10_cal = 16'b0000010011111011;
            15'd18038: log10_cal = 16'b0000010011111011;
            15'd18039: log10_cal = 16'b0000010011111011;
            15'd18040: log10_cal = 16'b0000010011111011;
            15'd18041: log10_cal = 16'b0000010011111011;
            15'd18042: log10_cal = 16'b0000010011111011;
            15'd18043: log10_cal = 16'b0000010011111011;
            15'd18044: log10_cal = 16'b0000010011111011;
            15'd18045: log10_cal = 16'b0000010011111011;
            15'd18046: log10_cal = 16'b0000010011111011;
            15'd18047: log10_cal = 16'b0000010011111100;
            15'd18048: log10_cal = 16'b0000010011111100;
            15'd18049: log10_cal = 16'b0000010011111100;
            15'd18050: log10_cal = 16'b0000010011111100;
            15'd18051: log10_cal = 16'b0000010011111100;
            15'd18052: log10_cal = 16'b0000010011111100;
            15'd18053: log10_cal = 16'b0000010011111100;
            15'd18054: log10_cal = 16'b0000010011111100;
            15'd18055: log10_cal = 16'b0000010011111100;
            15'd18056: log10_cal = 16'b0000010011111100;
            15'd18057: log10_cal = 16'b0000010011111100;
            15'd18058: log10_cal = 16'b0000010011111100;
            15'd18059: log10_cal = 16'b0000010011111100;
            15'd18060: log10_cal = 16'b0000010011111100;
            15'd18061: log10_cal = 16'b0000010011111100;
            15'd18062: log10_cal = 16'b0000010011111100;
            15'd18063: log10_cal = 16'b0000010011111100;
            15'd18064: log10_cal = 16'b0000010011111100;
            15'd18065: log10_cal = 16'b0000010011111100;
            15'd18066: log10_cal = 16'b0000010011111100;
            15'd18067: log10_cal = 16'b0000010011111100;
            15'd18068: log10_cal = 16'b0000010011111100;
            15'd18069: log10_cal = 16'b0000010011111100;
            15'd18070: log10_cal = 16'b0000010011111100;
            15'd18071: log10_cal = 16'b0000010011111100;
            15'd18072: log10_cal = 16'b0000010011111100;
            15'd18073: log10_cal = 16'b0000010011111100;
            15'd18074: log10_cal = 16'b0000010011111100;
            15'd18075: log10_cal = 16'b0000010011111100;
            15'd18076: log10_cal = 16'b0000010011111100;
            15'd18077: log10_cal = 16'b0000010011111100;
            15'd18078: log10_cal = 16'b0000010011111100;
            15'd18079: log10_cal = 16'b0000010011111100;
            15'd18080: log10_cal = 16'b0000010011111100;
            15'd18081: log10_cal = 16'b0000010011111100;
            15'd18082: log10_cal = 16'b0000010011111100;
            15'd18083: log10_cal = 16'b0000010011111100;
            15'd18084: log10_cal = 16'b0000010011111100;
            15'd18085: log10_cal = 16'b0000010011111100;
            15'd18086: log10_cal = 16'b0000010011111100;
            15'd18087: log10_cal = 16'b0000010011111100;
            15'd18088: log10_cal = 16'b0000010011111101;
            15'd18089: log10_cal = 16'b0000010011111101;
            15'd18090: log10_cal = 16'b0000010011111101;
            15'd18091: log10_cal = 16'b0000010011111101;
            15'd18092: log10_cal = 16'b0000010011111101;
            15'd18093: log10_cal = 16'b0000010011111101;
            15'd18094: log10_cal = 16'b0000010011111101;
            15'd18095: log10_cal = 16'b0000010011111101;
            15'd18096: log10_cal = 16'b0000010011111101;
            15'd18097: log10_cal = 16'b0000010011111101;
            15'd18098: log10_cal = 16'b0000010011111101;
            15'd18099: log10_cal = 16'b0000010011111101;
            15'd18100: log10_cal = 16'b0000010011111101;
            15'd18101: log10_cal = 16'b0000010011111101;
            15'd18102: log10_cal = 16'b0000010011111101;
            15'd18103: log10_cal = 16'b0000010011111101;
            15'd18104: log10_cal = 16'b0000010011111101;
            15'd18105: log10_cal = 16'b0000010011111101;
            15'd18106: log10_cal = 16'b0000010011111101;
            15'd18107: log10_cal = 16'b0000010011111101;
            15'd18108: log10_cal = 16'b0000010011111101;
            15'd18109: log10_cal = 16'b0000010011111101;
            15'd18110: log10_cal = 16'b0000010011111101;
            15'd18111: log10_cal = 16'b0000010011111101;
            15'd18112: log10_cal = 16'b0000010011111101;
            15'd18113: log10_cal = 16'b0000010011111101;
            15'd18114: log10_cal = 16'b0000010011111101;
            15'd18115: log10_cal = 16'b0000010011111101;
            15'd18116: log10_cal = 16'b0000010011111101;
            15'd18117: log10_cal = 16'b0000010011111101;
            15'd18118: log10_cal = 16'b0000010011111101;
            15'd18119: log10_cal = 16'b0000010011111101;
            15'd18120: log10_cal = 16'b0000010011111101;
            15'd18121: log10_cal = 16'b0000010011111101;
            15'd18122: log10_cal = 16'b0000010011111101;
            15'd18123: log10_cal = 16'b0000010011111101;
            15'd18124: log10_cal = 16'b0000010011111101;
            15'd18125: log10_cal = 16'b0000010011111101;
            15'd18126: log10_cal = 16'b0000010011111101;
            15'd18127: log10_cal = 16'b0000010011111101;
            15'd18128: log10_cal = 16'b0000010011111110;
            15'd18129: log10_cal = 16'b0000010011111110;
            15'd18130: log10_cal = 16'b0000010011111110;
            15'd18131: log10_cal = 16'b0000010011111110;
            15'd18132: log10_cal = 16'b0000010011111110;
            15'd18133: log10_cal = 16'b0000010011111110;
            15'd18134: log10_cal = 16'b0000010011111110;
            15'd18135: log10_cal = 16'b0000010011111110;
            15'd18136: log10_cal = 16'b0000010011111110;
            15'd18137: log10_cal = 16'b0000010011111110;
            15'd18138: log10_cal = 16'b0000010011111110;
            15'd18139: log10_cal = 16'b0000010011111110;
            15'd18140: log10_cal = 16'b0000010011111110;
            15'd18141: log10_cal = 16'b0000010011111110;
            15'd18142: log10_cal = 16'b0000010011111110;
            15'd18143: log10_cal = 16'b0000010011111110;
            15'd18144: log10_cal = 16'b0000010011111110;
            15'd18145: log10_cal = 16'b0000010011111110;
            15'd18146: log10_cal = 16'b0000010011111110;
            15'd18147: log10_cal = 16'b0000010011111110;
            15'd18148: log10_cal = 16'b0000010011111110;
            15'd18149: log10_cal = 16'b0000010011111110;
            15'd18150: log10_cal = 16'b0000010011111110;
            15'd18151: log10_cal = 16'b0000010011111110;
            15'd18152: log10_cal = 16'b0000010011111110;
            15'd18153: log10_cal = 16'b0000010011111110;
            15'd18154: log10_cal = 16'b0000010011111110;
            15'd18155: log10_cal = 16'b0000010011111110;
            15'd18156: log10_cal = 16'b0000010011111110;
            15'd18157: log10_cal = 16'b0000010011111110;
            15'd18158: log10_cal = 16'b0000010011111110;
            15'd18159: log10_cal = 16'b0000010011111110;
            15'd18160: log10_cal = 16'b0000010011111110;
            15'd18161: log10_cal = 16'b0000010011111110;
            15'd18162: log10_cal = 16'b0000010011111110;
            15'd18163: log10_cal = 16'b0000010011111110;
            15'd18164: log10_cal = 16'b0000010011111110;
            15'd18165: log10_cal = 16'b0000010011111110;
            15'd18166: log10_cal = 16'b0000010011111110;
            15'd18167: log10_cal = 16'b0000010011111110;
            15'd18168: log10_cal = 16'b0000010011111110;
            15'd18169: log10_cal = 16'b0000010011111111;
            15'd18170: log10_cal = 16'b0000010011111111;
            15'd18171: log10_cal = 16'b0000010011111111;
            15'd18172: log10_cal = 16'b0000010011111111;
            15'd18173: log10_cal = 16'b0000010011111111;
            15'd18174: log10_cal = 16'b0000010011111111;
            15'd18175: log10_cal = 16'b0000010011111111;
            15'd18176: log10_cal = 16'b0000010011111111;
            15'd18177: log10_cal = 16'b0000010011111111;
            15'd18178: log10_cal = 16'b0000010011111111;
            15'd18179: log10_cal = 16'b0000010011111111;
            15'd18180: log10_cal = 16'b0000010011111111;
            15'd18181: log10_cal = 16'b0000010011111111;
            15'd18182: log10_cal = 16'b0000010011111111;
            15'd18183: log10_cal = 16'b0000010011111111;
            15'd18184: log10_cal = 16'b0000010011111111;
            15'd18185: log10_cal = 16'b0000010011111111;
            15'd18186: log10_cal = 16'b0000010011111111;
            15'd18187: log10_cal = 16'b0000010011111111;
            15'd18188: log10_cal = 16'b0000010011111111;
            15'd18189: log10_cal = 16'b0000010011111111;
            15'd18190: log10_cal = 16'b0000010011111111;
            15'd18191: log10_cal = 16'b0000010011111111;
            15'd18192: log10_cal = 16'b0000010011111111;
            15'd18193: log10_cal = 16'b0000010011111111;
            15'd18194: log10_cal = 16'b0000010011111111;
            15'd18195: log10_cal = 16'b0000010011111111;
            15'd18196: log10_cal = 16'b0000010011111111;
            15'd18197: log10_cal = 16'b0000010011111111;
            15'd18198: log10_cal = 16'b0000010011111111;
            15'd18199: log10_cal = 16'b0000010011111111;
            15'd18200: log10_cal = 16'b0000010011111111;
            15'd18201: log10_cal = 16'b0000010011111111;
            15'd18202: log10_cal = 16'b0000010011111111;
            15'd18203: log10_cal = 16'b0000010011111111;
            15'd18204: log10_cal = 16'b0000010011111111;
            15'd18205: log10_cal = 16'b0000010011111111;
            15'd18206: log10_cal = 16'b0000010011111111;
            15'd18207: log10_cal = 16'b0000010011111111;
            15'd18208: log10_cal = 16'b0000010011111111;
            15'd18209: log10_cal = 16'b0000010011111111;
            15'd18210: log10_cal = 16'b0000010100000000;
            15'd18211: log10_cal = 16'b0000010100000000;
            15'd18212: log10_cal = 16'b0000010100000000;
            15'd18213: log10_cal = 16'b0000010100000000;
            15'd18214: log10_cal = 16'b0000010100000000;
            15'd18215: log10_cal = 16'b0000010100000000;
            15'd18216: log10_cal = 16'b0000010100000000;
            15'd18217: log10_cal = 16'b0000010100000000;
            15'd18218: log10_cal = 16'b0000010100000000;
            15'd18219: log10_cal = 16'b0000010100000000;
            15'd18220: log10_cal = 16'b0000010100000000;
            15'd18221: log10_cal = 16'b0000010100000000;
            15'd18222: log10_cal = 16'b0000010100000000;
            15'd18223: log10_cal = 16'b0000010100000000;
            15'd18224: log10_cal = 16'b0000010100000000;
            15'd18225: log10_cal = 16'b0000010100000000;
            15'd18226: log10_cal = 16'b0000010100000000;
            15'd18227: log10_cal = 16'b0000010100000000;
            15'd18228: log10_cal = 16'b0000010100000000;
            15'd18229: log10_cal = 16'b0000010100000000;
            15'd18230: log10_cal = 16'b0000010100000000;
            15'd18231: log10_cal = 16'b0000010100000000;
            15'd18232: log10_cal = 16'b0000010100000000;
            15'd18233: log10_cal = 16'b0000010100000000;
            15'd18234: log10_cal = 16'b0000010100000000;
            15'd18235: log10_cal = 16'b0000010100000000;
            15'd18236: log10_cal = 16'b0000010100000000;
            15'd18237: log10_cal = 16'b0000010100000000;
            15'd18238: log10_cal = 16'b0000010100000000;
            15'd18239: log10_cal = 16'b0000010100000000;
            15'd18240: log10_cal = 16'b0000010100000000;
            15'd18241: log10_cal = 16'b0000010100000000;
            15'd18242: log10_cal = 16'b0000010100000000;
            15'd18243: log10_cal = 16'b0000010100000000;
            15'd18244: log10_cal = 16'b0000010100000000;
            15'd18245: log10_cal = 16'b0000010100000000;
            15'd18246: log10_cal = 16'b0000010100000000;
            15'd18247: log10_cal = 16'b0000010100000000;
            15'd18248: log10_cal = 16'b0000010100000000;
            15'd18249: log10_cal = 16'b0000010100000000;
            15'd18250: log10_cal = 16'b0000010100000000;
            15'd18251: log10_cal = 16'b0000010100000001;
            15'd18252: log10_cal = 16'b0000010100000001;
            15'd18253: log10_cal = 16'b0000010100000001;
            15'd18254: log10_cal = 16'b0000010100000001;
            15'd18255: log10_cal = 16'b0000010100000001;
            15'd18256: log10_cal = 16'b0000010100000001;
            15'd18257: log10_cal = 16'b0000010100000001;
            15'd18258: log10_cal = 16'b0000010100000001;
            15'd18259: log10_cal = 16'b0000010100000001;
            15'd18260: log10_cal = 16'b0000010100000001;
            15'd18261: log10_cal = 16'b0000010100000001;
            15'd18262: log10_cal = 16'b0000010100000001;
            15'd18263: log10_cal = 16'b0000010100000001;
            15'd18264: log10_cal = 16'b0000010100000001;
            15'd18265: log10_cal = 16'b0000010100000001;
            15'd18266: log10_cal = 16'b0000010100000001;
            15'd18267: log10_cal = 16'b0000010100000001;
            15'd18268: log10_cal = 16'b0000010100000001;
            15'd18269: log10_cal = 16'b0000010100000001;
            15'd18270: log10_cal = 16'b0000010100000001;
            15'd18271: log10_cal = 16'b0000010100000001;
            15'd18272: log10_cal = 16'b0000010100000001;
            15'd18273: log10_cal = 16'b0000010100000001;
            15'd18274: log10_cal = 16'b0000010100000001;
            15'd18275: log10_cal = 16'b0000010100000001;
            15'd18276: log10_cal = 16'b0000010100000001;
            15'd18277: log10_cal = 16'b0000010100000001;
            15'd18278: log10_cal = 16'b0000010100000001;
            15'd18279: log10_cal = 16'b0000010100000001;
            15'd18280: log10_cal = 16'b0000010100000001;
            15'd18281: log10_cal = 16'b0000010100000001;
            15'd18282: log10_cal = 16'b0000010100000001;
            15'd18283: log10_cal = 16'b0000010100000001;
            15'd18284: log10_cal = 16'b0000010100000001;
            15'd18285: log10_cal = 16'b0000010100000001;
            15'd18286: log10_cal = 16'b0000010100000001;
            15'd18287: log10_cal = 16'b0000010100000001;
            15'd18288: log10_cal = 16'b0000010100000001;
            15'd18289: log10_cal = 16'b0000010100000001;
            15'd18290: log10_cal = 16'b0000010100000001;
            15'd18291: log10_cal = 16'b0000010100000001;
            15'd18292: log10_cal = 16'b0000010100000010;
            15'd18293: log10_cal = 16'b0000010100000010;
            15'd18294: log10_cal = 16'b0000010100000010;
            15'd18295: log10_cal = 16'b0000010100000010;
            15'd18296: log10_cal = 16'b0000010100000010;
            15'd18297: log10_cal = 16'b0000010100000010;
            15'd18298: log10_cal = 16'b0000010100000010;
            15'd18299: log10_cal = 16'b0000010100000010;
            15'd18300: log10_cal = 16'b0000010100000010;
            15'd18301: log10_cal = 16'b0000010100000010;
            15'd18302: log10_cal = 16'b0000010100000010;
            15'd18303: log10_cal = 16'b0000010100000010;
            15'd18304: log10_cal = 16'b0000010100000010;
            15'd18305: log10_cal = 16'b0000010100000010;
            15'd18306: log10_cal = 16'b0000010100000010;
            15'd18307: log10_cal = 16'b0000010100000010;
            15'd18308: log10_cal = 16'b0000010100000010;
            15'd18309: log10_cal = 16'b0000010100000010;
            15'd18310: log10_cal = 16'b0000010100000010;
            15'd18311: log10_cal = 16'b0000010100000010;
            15'd18312: log10_cal = 16'b0000010100000010;
            15'd18313: log10_cal = 16'b0000010100000010;
            15'd18314: log10_cal = 16'b0000010100000010;
            15'd18315: log10_cal = 16'b0000010100000010;
            15'd18316: log10_cal = 16'b0000010100000010;
            15'd18317: log10_cal = 16'b0000010100000010;
            15'd18318: log10_cal = 16'b0000010100000010;
            15'd18319: log10_cal = 16'b0000010100000010;
            15'd18320: log10_cal = 16'b0000010100000010;
            15'd18321: log10_cal = 16'b0000010100000010;
            15'd18322: log10_cal = 16'b0000010100000010;
            15'd18323: log10_cal = 16'b0000010100000010;
            15'd18324: log10_cal = 16'b0000010100000010;
            15'd18325: log10_cal = 16'b0000010100000010;
            15'd18326: log10_cal = 16'b0000010100000010;
            15'd18327: log10_cal = 16'b0000010100000010;
            15'd18328: log10_cal = 16'b0000010100000010;
            15'd18329: log10_cal = 16'b0000010100000010;
            15'd18330: log10_cal = 16'b0000010100000010;
            15'd18331: log10_cal = 16'b0000010100000010;
            15'd18332: log10_cal = 16'b0000010100000010;
            15'd18333: log10_cal = 16'b0000010100000011;
            15'd18334: log10_cal = 16'b0000010100000011;
            15'd18335: log10_cal = 16'b0000010100000011;
            15'd18336: log10_cal = 16'b0000010100000011;
            15'd18337: log10_cal = 16'b0000010100000011;
            15'd18338: log10_cal = 16'b0000010100000011;
            15'd18339: log10_cal = 16'b0000010100000011;
            15'd18340: log10_cal = 16'b0000010100000011;
            15'd18341: log10_cal = 16'b0000010100000011;
            15'd18342: log10_cal = 16'b0000010100000011;
            15'd18343: log10_cal = 16'b0000010100000011;
            15'd18344: log10_cal = 16'b0000010100000011;
            15'd18345: log10_cal = 16'b0000010100000011;
            15'd18346: log10_cal = 16'b0000010100000011;
            15'd18347: log10_cal = 16'b0000010100000011;
            15'd18348: log10_cal = 16'b0000010100000011;
            15'd18349: log10_cal = 16'b0000010100000011;
            15'd18350: log10_cal = 16'b0000010100000011;
            15'd18351: log10_cal = 16'b0000010100000011;
            15'd18352: log10_cal = 16'b0000010100000011;
            15'd18353: log10_cal = 16'b0000010100000011;
            15'd18354: log10_cal = 16'b0000010100000011;
            15'd18355: log10_cal = 16'b0000010100000011;
            15'd18356: log10_cal = 16'b0000010100000011;
            15'd18357: log10_cal = 16'b0000010100000011;
            15'd18358: log10_cal = 16'b0000010100000011;
            15'd18359: log10_cal = 16'b0000010100000011;
            15'd18360: log10_cal = 16'b0000010100000011;
            15'd18361: log10_cal = 16'b0000010100000011;
            15'd18362: log10_cal = 16'b0000010100000011;
            15'd18363: log10_cal = 16'b0000010100000011;
            15'd18364: log10_cal = 16'b0000010100000011;
            15'd18365: log10_cal = 16'b0000010100000011;
            15'd18366: log10_cal = 16'b0000010100000011;
            15'd18367: log10_cal = 16'b0000010100000011;
            15'd18368: log10_cal = 16'b0000010100000011;
            15'd18369: log10_cal = 16'b0000010100000011;
            15'd18370: log10_cal = 16'b0000010100000011;
            15'd18371: log10_cal = 16'b0000010100000011;
            15'd18372: log10_cal = 16'b0000010100000011;
            15'd18373: log10_cal = 16'b0000010100000011;
            15'd18374: log10_cal = 16'b0000010100000011;
            15'd18375: log10_cal = 16'b0000010100000100;
            15'd18376: log10_cal = 16'b0000010100000100;
            15'd18377: log10_cal = 16'b0000010100000100;
            15'd18378: log10_cal = 16'b0000010100000100;
            15'd18379: log10_cal = 16'b0000010100000100;
            15'd18380: log10_cal = 16'b0000010100000100;
            15'd18381: log10_cal = 16'b0000010100000100;
            15'd18382: log10_cal = 16'b0000010100000100;
            15'd18383: log10_cal = 16'b0000010100000100;
            15'd18384: log10_cal = 16'b0000010100000100;
            15'd18385: log10_cal = 16'b0000010100000100;
            15'd18386: log10_cal = 16'b0000010100000100;
            15'd18387: log10_cal = 16'b0000010100000100;
            15'd18388: log10_cal = 16'b0000010100000100;
            15'd18389: log10_cal = 16'b0000010100000100;
            15'd18390: log10_cal = 16'b0000010100000100;
            15'd18391: log10_cal = 16'b0000010100000100;
            15'd18392: log10_cal = 16'b0000010100000100;
            15'd18393: log10_cal = 16'b0000010100000100;
            15'd18394: log10_cal = 16'b0000010100000100;
            15'd18395: log10_cal = 16'b0000010100000100;
            15'd18396: log10_cal = 16'b0000010100000100;
            15'd18397: log10_cal = 16'b0000010100000100;
            15'd18398: log10_cal = 16'b0000010100000100;
            15'd18399: log10_cal = 16'b0000010100000100;
            15'd18400: log10_cal = 16'b0000010100000100;
            15'd18401: log10_cal = 16'b0000010100000100;
            15'd18402: log10_cal = 16'b0000010100000100;
            15'd18403: log10_cal = 16'b0000010100000100;
            15'd18404: log10_cal = 16'b0000010100000100;
            15'd18405: log10_cal = 16'b0000010100000100;
            15'd18406: log10_cal = 16'b0000010100000100;
            15'd18407: log10_cal = 16'b0000010100000100;
            15'd18408: log10_cal = 16'b0000010100000100;
            15'd18409: log10_cal = 16'b0000010100000100;
            15'd18410: log10_cal = 16'b0000010100000100;
            15'd18411: log10_cal = 16'b0000010100000100;
            15'd18412: log10_cal = 16'b0000010100000100;
            15'd18413: log10_cal = 16'b0000010100000100;
            15'd18414: log10_cal = 16'b0000010100000100;
            15'd18415: log10_cal = 16'b0000010100000100;
            15'd18416: log10_cal = 16'b0000010100000101;
            15'd18417: log10_cal = 16'b0000010100000101;
            15'd18418: log10_cal = 16'b0000010100000101;
            15'd18419: log10_cal = 16'b0000010100000101;
            15'd18420: log10_cal = 16'b0000010100000101;
            15'd18421: log10_cal = 16'b0000010100000101;
            15'd18422: log10_cal = 16'b0000010100000101;
            15'd18423: log10_cal = 16'b0000010100000101;
            15'd18424: log10_cal = 16'b0000010100000101;
            15'd18425: log10_cal = 16'b0000010100000101;
            15'd18426: log10_cal = 16'b0000010100000101;
            15'd18427: log10_cal = 16'b0000010100000101;
            15'd18428: log10_cal = 16'b0000010100000101;
            15'd18429: log10_cal = 16'b0000010100000101;
            15'd18430: log10_cal = 16'b0000010100000101;
            15'd18431: log10_cal = 16'b0000010100000101;
            15'd18432: log10_cal = 16'b0000010100000101;
            15'd18433: log10_cal = 16'b0000010100000101;
            15'd18434: log10_cal = 16'b0000010100000101;
            15'd18435: log10_cal = 16'b0000010100000101;
            15'd18436: log10_cal = 16'b0000010100000101;
            15'd18437: log10_cal = 16'b0000010100000101;
            15'd18438: log10_cal = 16'b0000010100000101;
            15'd18439: log10_cal = 16'b0000010100000101;
            15'd18440: log10_cal = 16'b0000010100000101;
            15'd18441: log10_cal = 16'b0000010100000101;
            15'd18442: log10_cal = 16'b0000010100000101;
            15'd18443: log10_cal = 16'b0000010100000101;
            15'd18444: log10_cal = 16'b0000010100000101;
            15'd18445: log10_cal = 16'b0000010100000101;
            15'd18446: log10_cal = 16'b0000010100000101;
            15'd18447: log10_cal = 16'b0000010100000101;
            15'd18448: log10_cal = 16'b0000010100000101;
            15'd18449: log10_cal = 16'b0000010100000101;
            15'd18450: log10_cal = 16'b0000010100000101;
            15'd18451: log10_cal = 16'b0000010100000101;
            15'd18452: log10_cal = 16'b0000010100000101;
            15'd18453: log10_cal = 16'b0000010100000101;
            15'd18454: log10_cal = 16'b0000010100000101;
            15'd18455: log10_cal = 16'b0000010100000101;
            15'd18456: log10_cal = 16'b0000010100000101;
            15'd18457: log10_cal = 16'b0000010100000110;
            15'd18458: log10_cal = 16'b0000010100000110;
            15'd18459: log10_cal = 16'b0000010100000110;
            15'd18460: log10_cal = 16'b0000010100000110;
            15'd18461: log10_cal = 16'b0000010100000110;
            15'd18462: log10_cal = 16'b0000010100000110;
            15'd18463: log10_cal = 16'b0000010100000110;
            15'd18464: log10_cal = 16'b0000010100000110;
            15'd18465: log10_cal = 16'b0000010100000110;
            15'd18466: log10_cal = 16'b0000010100000110;
            15'd18467: log10_cal = 16'b0000010100000110;
            15'd18468: log10_cal = 16'b0000010100000110;
            15'd18469: log10_cal = 16'b0000010100000110;
            15'd18470: log10_cal = 16'b0000010100000110;
            15'd18471: log10_cal = 16'b0000010100000110;
            15'd18472: log10_cal = 16'b0000010100000110;
            15'd18473: log10_cal = 16'b0000010100000110;
            15'd18474: log10_cal = 16'b0000010100000110;
            15'd18475: log10_cal = 16'b0000010100000110;
            15'd18476: log10_cal = 16'b0000010100000110;
            15'd18477: log10_cal = 16'b0000010100000110;
            15'd18478: log10_cal = 16'b0000010100000110;
            15'd18479: log10_cal = 16'b0000010100000110;
            15'd18480: log10_cal = 16'b0000010100000110;
            15'd18481: log10_cal = 16'b0000010100000110;
            15'd18482: log10_cal = 16'b0000010100000110;
            15'd18483: log10_cal = 16'b0000010100000110;
            15'd18484: log10_cal = 16'b0000010100000110;
            15'd18485: log10_cal = 16'b0000010100000110;
            15'd18486: log10_cal = 16'b0000010100000110;
            15'd18487: log10_cal = 16'b0000010100000110;
            15'd18488: log10_cal = 16'b0000010100000110;
            15'd18489: log10_cal = 16'b0000010100000110;
            15'd18490: log10_cal = 16'b0000010100000110;
            15'd18491: log10_cal = 16'b0000010100000110;
            15'd18492: log10_cal = 16'b0000010100000110;
            15'd18493: log10_cal = 16'b0000010100000110;
            15'd18494: log10_cal = 16'b0000010100000110;
            15'd18495: log10_cal = 16'b0000010100000110;
            15'd18496: log10_cal = 16'b0000010100000110;
            15'd18497: log10_cal = 16'b0000010100000110;
            15'd18498: log10_cal = 16'b0000010100000110;
            15'd18499: log10_cal = 16'b0000010100000111;
            15'd18500: log10_cal = 16'b0000010100000111;
            15'd18501: log10_cal = 16'b0000010100000111;
            15'd18502: log10_cal = 16'b0000010100000111;
            15'd18503: log10_cal = 16'b0000010100000111;
            15'd18504: log10_cal = 16'b0000010100000111;
            15'd18505: log10_cal = 16'b0000010100000111;
            15'd18506: log10_cal = 16'b0000010100000111;
            15'd18507: log10_cal = 16'b0000010100000111;
            15'd18508: log10_cal = 16'b0000010100000111;
            15'd18509: log10_cal = 16'b0000010100000111;
            15'd18510: log10_cal = 16'b0000010100000111;
            15'd18511: log10_cal = 16'b0000010100000111;
            15'd18512: log10_cal = 16'b0000010100000111;
            15'd18513: log10_cal = 16'b0000010100000111;
            15'd18514: log10_cal = 16'b0000010100000111;
            15'd18515: log10_cal = 16'b0000010100000111;
            15'd18516: log10_cal = 16'b0000010100000111;
            15'd18517: log10_cal = 16'b0000010100000111;
            15'd18518: log10_cal = 16'b0000010100000111;
            15'd18519: log10_cal = 16'b0000010100000111;
            15'd18520: log10_cal = 16'b0000010100000111;
            15'd18521: log10_cal = 16'b0000010100000111;
            15'd18522: log10_cal = 16'b0000010100000111;
            15'd18523: log10_cal = 16'b0000010100000111;
            15'd18524: log10_cal = 16'b0000010100000111;
            15'd18525: log10_cal = 16'b0000010100000111;
            15'd18526: log10_cal = 16'b0000010100000111;
            15'd18527: log10_cal = 16'b0000010100000111;
            15'd18528: log10_cal = 16'b0000010100000111;
            15'd18529: log10_cal = 16'b0000010100000111;
            15'd18530: log10_cal = 16'b0000010100000111;
            15'd18531: log10_cal = 16'b0000010100000111;
            15'd18532: log10_cal = 16'b0000010100000111;
            15'd18533: log10_cal = 16'b0000010100000111;
            15'd18534: log10_cal = 16'b0000010100000111;
            15'd18535: log10_cal = 16'b0000010100000111;
            15'd18536: log10_cal = 16'b0000010100000111;
            15'd18537: log10_cal = 16'b0000010100000111;
            15'd18538: log10_cal = 16'b0000010100000111;
            15'd18539: log10_cal = 16'b0000010100000111;
            15'd18540: log10_cal = 16'b0000010100000111;
            15'd18541: log10_cal = 16'b0000010100001000;
            15'd18542: log10_cal = 16'b0000010100001000;
            15'd18543: log10_cal = 16'b0000010100001000;
            15'd18544: log10_cal = 16'b0000010100001000;
            15'd18545: log10_cal = 16'b0000010100001000;
            15'd18546: log10_cal = 16'b0000010100001000;
            15'd18547: log10_cal = 16'b0000010100001000;
            15'd18548: log10_cal = 16'b0000010100001000;
            15'd18549: log10_cal = 16'b0000010100001000;
            15'd18550: log10_cal = 16'b0000010100001000;
            15'd18551: log10_cal = 16'b0000010100001000;
            15'd18552: log10_cal = 16'b0000010100001000;
            15'd18553: log10_cal = 16'b0000010100001000;
            15'd18554: log10_cal = 16'b0000010100001000;
            15'd18555: log10_cal = 16'b0000010100001000;
            15'd18556: log10_cal = 16'b0000010100001000;
            15'd18557: log10_cal = 16'b0000010100001000;
            15'd18558: log10_cal = 16'b0000010100001000;
            15'd18559: log10_cal = 16'b0000010100001000;
            15'd18560: log10_cal = 16'b0000010100001000;
            15'd18561: log10_cal = 16'b0000010100001000;
            15'd18562: log10_cal = 16'b0000010100001000;
            15'd18563: log10_cal = 16'b0000010100001000;
            15'd18564: log10_cal = 16'b0000010100001000;
            15'd18565: log10_cal = 16'b0000010100001000;
            15'd18566: log10_cal = 16'b0000010100001000;
            15'd18567: log10_cal = 16'b0000010100001000;
            15'd18568: log10_cal = 16'b0000010100001000;
            15'd18569: log10_cal = 16'b0000010100001000;
            15'd18570: log10_cal = 16'b0000010100001000;
            15'd18571: log10_cal = 16'b0000010100001000;
            15'd18572: log10_cal = 16'b0000010100001000;
            15'd18573: log10_cal = 16'b0000010100001000;
            15'd18574: log10_cal = 16'b0000010100001000;
            15'd18575: log10_cal = 16'b0000010100001000;
            15'd18576: log10_cal = 16'b0000010100001000;
            15'd18577: log10_cal = 16'b0000010100001000;
            15'd18578: log10_cal = 16'b0000010100001000;
            15'd18579: log10_cal = 16'b0000010100001000;
            15'd18580: log10_cal = 16'b0000010100001000;
            15'd18581: log10_cal = 16'b0000010100001000;
            15'd18582: log10_cal = 16'b0000010100001001;
            15'd18583: log10_cal = 16'b0000010100001001;
            15'd18584: log10_cal = 16'b0000010100001001;
            15'd18585: log10_cal = 16'b0000010100001001;
            15'd18586: log10_cal = 16'b0000010100001001;
            15'd18587: log10_cal = 16'b0000010100001001;
            15'd18588: log10_cal = 16'b0000010100001001;
            15'd18589: log10_cal = 16'b0000010100001001;
            15'd18590: log10_cal = 16'b0000010100001001;
            15'd18591: log10_cal = 16'b0000010100001001;
            15'd18592: log10_cal = 16'b0000010100001001;
            15'd18593: log10_cal = 16'b0000010100001001;
            15'd18594: log10_cal = 16'b0000010100001001;
            15'd18595: log10_cal = 16'b0000010100001001;
            15'd18596: log10_cal = 16'b0000010100001001;
            15'd18597: log10_cal = 16'b0000010100001001;
            15'd18598: log10_cal = 16'b0000010100001001;
            15'd18599: log10_cal = 16'b0000010100001001;
            15'd18600: log10_cal = 16'b0000010100001001;
            15'd18601: log10_cal = 16'b0000010100001001;
            15'd18602: log10_cal = 16'b0000010100001001;
            15'd18603: log10_cal = 16'b0000010100001001;
            15'd18604: log10_cal = 16'b0000010100001001;
            15'd18605: log10_cal = 16'b0000010100001001;
            15'd18606: log10_cal = 16'b0000010100001001;
            15'd18607: log10_cal = 16'b0000010100001001;
            15'd18608: log10_cal = 16'b0000010100001001;
            15'd18609: log10_cal = 16'b0000010100001001;
            15'd18610: log10_cal = 16'b0000010100001001;
            15'd18611: log10_cal = 16'b0000010100001001;
            15'd18612: log10_cal = 16'b0000010100001001;
            15'd18613: log10_cal = 16'b0000010100001001;
            15'd18614: log10_cal = 16'b0000010100001001;
            15'd18615: log10_cal = 16'b0000010100001001;
            15'd18616: log10_cal = 16'b0000010100001001;
            15'd18617: log10_cal = 16'b0000010100001001;
            15'd18618: log10_cal = 16'b0000010100001001;
            15'd18619: log10_cal = 16'b0000010100001001;
            15'd18620: log10_cal = 16'b0000010100001001;
            15'd18621: log10_cal = 16'b0000010100001001;
            15'd18622: log10_cal = 16'b0000010100001001;
            15'd18623: log10_cal = 16'b0000010100001001;
            15'd18624: log10_cal = 16'b0000010100001010;
            15'd18625: log10_cal = 16'b0000010100001010;
            15'd18626: log10_cal = 16'b0000010100001010;
            15'd18627: log10_cal = 16'b0000010100001010;
            15'd18628: log10_cal = 16'b0000010100001010;
            15'd18629: log10_cal = 16'b0000010100001010;
            15'd18630: log10_cal = 16'b0000010100001010;
            15'd18631: log10_cal = 16'b0000010100001010;
            15'd18632: log10_cal = 16'b0000010100001010;
            15'd18633: log10_cal = 16'b0000010100001010;
            15'd18634: log10_cal = 16'b0000010100001010;
            15'd18635: log10_cal = 16'b0000010100001010;
            15'd18636: log10_cal = 16'b0000010100001010;
            15'd18637: log10_cal = 16'b0000010100001010;
            15'd18638: log10_cal = 16'b0000010100001010;
            15'd18639: log10_cal = 16'b0000010100001010;
            15'd18640: log10_cal = 16'b0000010100001010;
            15'd18641: log10_cal = 16'b0000010100001010;
            15'd18642: log10_cal = 16'b0000010100001010;
            15'd18643: log10_cal = 16'b0000010100001010;
            15'd18644: log10_cal = 16'b0000010100001010;
            15'd18645: log10_cal = 16'b0000010100001010;
            15'd18646: log10_cal = 16'b0000010100001010;
            15'd18647: log10_cal = 16'b0000010100001010;
            15'd18648: log10_cal = 16'b0000010100001010;
            15'd18649: log10_cal = 16'b0000010100001010;
            15'd18650: log10_cal = 16'b0000010100001010;
            15'd18651: log10_cal = 16'b0000010100001010;
            15'd18652: log10_cal = 16'b0000010100001010;
            15'd18653: log10_cal = 16'b0000010100001010;
            15'd18654: log10_cal = 16'b0000010100001010;
            15'd18655: log10_cal = 16'b0000010100001010;
            15'd18656: log10_cal = 16'b0000010100001010;
            15'd18657: log10_cal = 16'b0000010100001010;
            15'd18658: log10_cal = 16'b0000010100001010;
            15'd18659: log10_cal = 16'b0000010100001010;
            15'd18660: log10_cal = 16'b0000010100001010;
            15'd18661: log10_cal = 16'b0000010100001010;
            15'd18662: log10_cal = 16'b0000010100001010;
            15'd18663: log10_cal = 16'b0000010100001010;
            15'd18664: log10_cal = 16'b0000010100001010;
            15'd18665: log10_cal = 16'b0000010100001010;
            15'd18666: log10_cal = 16'b0000010100001011;
            15'd18667: log10_cal = 16'b0000010100001011;
            15'd18668: log10_cal = 16'b0000010100001011;
            15'd18669: log10_cal = 16'b0000010100001011;
            15'd18670: log10_cal = 16'b0000010100001011;
            15'd18671: log10_cal = 16'b0000010100001011;
            15'd18672: log10_cal = 16'b0000010100001011;
            15'd18673: log10_cal = 16'b0000010100001011;
            15'd18674: log10_cal = 16'b0000010100001011;
            15'd18675: log10_cal = 16'b0000010100001011;
            15'd18676: log10_cal = 16'b0000010100001011;
            15'd18677: log10_cal = 16'b0000010100001011;
            15'd18678: log10_cal = 16'b0000010100001011;
            15'd18679: log10_cal = 16'b0000010100001011;
            15'd18680: log10_cal = 16'b0000010100001011;
            15'd18681: log10_cal = 16'b0000010100001011;
            15'd18682: log10_cal = 16'b0000010100001011;
            15'd18683: log10_cal = 16'b0000010100001011;
            15'd18684: log10_cal = 16'b0000010100001011;
            15'd18685: log10_cal = 16'b0000010100001011;
            15'd18686: log10_cal = 16'b0000010100001011;
            15'd18687: log10_cal = 16'b0000010100001011;
            15'd18688: log10_cal = 16'b0000010100001011;
            15'd18689: log10_cal = 16'b0000010100001011;
            15'd18690: log10_cal = 16'b0000010100001011;
            15'd18691: log10_cal = 16'b0000010100001011;
            15'd18692: log10_cal = 16'b0000010100001011;
            15'd18693: log10_cal = 16'b0000010100001011;
            15'd18694: log10_cal = 16'b0000010100001011;
            15'd18695: log10_cal = 16'b0000010100001011;
            15'd18696: log10_cal = 16'b0000010100001011;
            15'd18697: log10_cal = 16'b0000010100001011;
            15'd18698: log10_cal = 16'b0000010100001011;
            15'd18699: log10_cal = 16'b0000010100001011;
            15'd18700: log10_cal = 16'b0000010100001011;
            15'd18701: log10_cal = 16'b0000010100001011;
            15'd18702: log10_cal = 16'b0000010100001011;
            15'd18703: log10_cal = 16'b0000010100001011;
            15'd18704: log10_cal = 16'b0000010100001011;
            15'd18705: log10_cal = 16'b0000010100001011;
            15'd18706: log10_cal = 16'b0000010100001011;
            15'd18707: log10_cal = 16'b0000010100001011;
            15'd18708: log10_cal = 16'b0000010100001100;
            15'd18709: log10_cal = 16'b0000010100001100;
            15'd18710: log10_cal = 16'b0000010100001100;
            15'd18711: log10_cal = 16'b0000010100001100;
            15'd18712: log10_cal = 16'b0000010100001100;
            15'd18713: log10_cal = 16'b0000010100001100;
            15'd18714: log10_cal = 16'b0000010100001100;
            15'd18715: log10_cal = 16'b0000010100001100;
            15'd18716: log10_cal = 16'b0000010100001100;
            15'd18717: log10_cal = 16'b0000010100001100;
            15'd18718: log10_cal = 16'b0000010100001100;
            15'd18719: log10_cal = 16'b0000010100001100;
            15'd18720: log10_cal = 16'b0000010100001100;
            15'd18721: log10_cal = 16'b0000010100001100;
            15'd18722: log10_cal = 16'b0000010100001100;
            15'd18723: log10_cal = 16'b0000010100001100;
            15'd18724: log10_cal = 16'b0000010100001100;
            15'd18725: log10_cal = 16'b0000010100001100;
            15'd18726: log10_cal = 16'b0000010100001100;
            15'd18727: log10_cal = 16'b0000010100001100;
            15'd18728: log10_cal = 16'b0000010100001100;
            15'd18729: log10_cal = 16'b0000010100001100;
            15'd18730: log10_cal = 16'b0000010100001100;
            15'd18731: log10_cal = 16'b0000010100001100;
            15'd18732: log10_cal = 16'b0000010100001100;
            15'd18733: log10_cal = 16'b0000010100001100;
            15'd18734: log10_cal = 16'b0000010100001100;
            15'd18735: log10_cal = 16'b0000010100001100;
            15'd18736: log10_cal = 16'b0000010100001100;
            15'd18737: log10_cal = 16'b0000010100001100;
            15'd18738: log10_cal = 16'b0000010100001100;
            15'd18739: log10_cal = 16'b0000010100001100;
            15'd18740: log10_cal = 16'b0000010100001100;
            15'd18741: log10_cal = 16'b0000010100001100;
            15'd18742: log10_cal = 16'b0000010100001100;
            15'd18743: log10_cal = 16'b0000010100001100;
            15'd18744: log10_cal = 16'b0000010100001100;
            15'd18745: log10_cal = 16'b0000010100001100;
            15'd18746: log10_cal = 16'b0000010100001100;
            15'd18747: log10_cal = 16'b0000010100001100;
            15'd18748: log10_cal = 16'b0000010100001100;
            15'd18749: log10_cal = 16'b0000010100001100;
            15'd18750: log10_cal = 16'b0000010100001101;
            15'd18751: log10_cal = 16'b0000010100001101;
            15'd18752: log10_cal = 16'b0000010100001101;
            15'd18753: log10_cal = 16'b0000010100001101;
            15'd18754: log10_cal = 16'b0000010100001101;
            15'd18755: log10_cal = 16'b0000010100001101;
            15'd18756: log10_cal = 16'b0000010100001101;
            15'd18757: log10_cal = 16'b0000010100001101;
            15'd18758: log10_cal = 16'b0000010100001101;
            15'd18759: log10_cal = 16'b0000010100001101;
            15'd18760: log10_cal = 16'b0000010100001101;
            15'd18761: log10_cal = 16'b0000010100001101;
            15'd18762: log10_cal = 16'b0000010100001101;
            15'd18763: log10_cal = 16'b0000010100001101;
            15'd18764: log10_cal = 16'b0000010100001101;
            15'd18765: log10_cal = 16'b0000010100001101;
            15'd18766: log10_cal = 16'b0000010100001101;
            15'd18767: log10_cal = 16'b0000010100001101;
            15'd18768: log10_cal = 16'b0000010100001101;
            15'd18769: log10_cal = 16'b0000010100001101;
            15'd18770: log10_cal = 16'b0000010100001101;
            15'd18771: log10_cal = 16'b0000010100001101;
            15'd18772: log10_cal = 16'b0000010100001101;
            15'd18773: log10_cal = 16'b0000010100001101;
            15'd18774: log10_cal = 16'b0000010100001101;
            15'd18775: log10_cal = 16'b0000010100001101;
            15'd18776: log10_cal = 16'b0000010100001101;
            15'd18777: log10_cal = 16'b0000010100001101;
            15'd18778: log10_cal = 16'b0000010100001101;
            15'd18779: log10_cal = 16'b0000010100001101;
            15'd18780: log10_cal = 16'b0000010100001101;
            15'd18781: log10_cal = 16'b0000010100001101;
            15'd18782: log10_cal = 16'b0000010100001101;
            15'd18783: log10_cal = 16'b0000010100001101;
            15'd18784: log10_cal = 16'b0000010100001101;
            15'd18785: log10_cal = 16'b0000010100001101;
            15'd18786: log10_cal = 16'b0000010100001101;
            15'd18787: log10_cal = 16'b0000010100001101;
            15'd18788: log10_cal = 16'b0000010100001101;
            15'd18789: log10_cal = 16'b0000010100001101;
            15'd18790: log10_cal = 16'b0000010100001101;
            15'd18791: log10_cal = 16'b0000010100001101;
            15'd18792: log10_cal = 16'b0000010100001110;
            15'd18793: log10_cal = 16'b0000010100001110;
            15'd18794: log10_cal = 16'b0000010100001110;
            15'd18795: log10_cal = 16'b0000010100001110;
            15'd18796: log10_cal = 16'b0000010100001110;
            15'd18797: log10_cal = 16'b0000010100001110;
            15'd18798: log10_cal = 16'b0000010100001110;
            15'd18799: log10_cal = 16'b0000010100001110;
            15'd18800: log10_cal = 16'b0000010100001110;
            15'd18801: log10_cal = 16'b0000010100001110;
            15'd18802: log10_cal = 16'b0000010100001110;
            15'd18803: log10_cal = 16'b0000010100001110;
            15'd18804: log10_cal = 16'b0000010100001110;
            15'd18805: log10_cal = 16'b0000010100001110;
            15'd18806: log10_cal = 16'b0000010100001110;
            15'd18807: log10_cal = 16'b0000010100001110;
            15'd18808: log10_cal = 16'b0000010100001110;
            15'd18809: log10_cal = 16'b0000010100001110;
            15'd18810: log10_cal = 16'b0000010100001110;
            15'd18811: log10_cal = 16'b0000010100001110;
            15'd18812: log10_cal = 16'b0000010100001110;
            15'd18813: log10_cal = 16'b0000010100001110;
            15'd18814: log10_cal = 16'b0000010100001110;
            15'd18815: log10_cal = 16'b0000010100001110;
            15'd18816: log10_cal = 16'b0000010100001110;
            15'd18817: log10_cal = 16'b0000010100001110;
            15'd18818: log10_cal = 16'b0000010100001110;
            15'd18819: log10_cal = 16'b0000010100001110;
            15'd18820: log10_cal = 16'b0000010100001110;
            15'd18821: log10_cal = 16'b0000010100001110;
            15'd18822: log10_cal = 16'b0000010100001110;
            15'd18823: log10_cal = 16'b0000010100001110;
            15'd18824: log10_cal = 16'b0000010100001110;
            15'd18825: log10_cal = 16'b0000010100001110;
            15'd18826: log10_cal = 16'b0000010100001110;
            15'd18827: log10_cal = 16'b0000010100001110;
            15'd18828: log10_cal = 16'b0000010100001110;
            15'd18829: log10_cal = 16'b0000010100001110;
            15'd18830: log10_cal = 16'b0000010100001110;
            15'd18831: log10_cal = 16'b0000010100001110;
            15'd18832: log10_cal = 16'b0000010100001110;
            15'd18833: log10_cal = 16'b0000010100001110;
            15'd18834: log10_cal = 16'b0000010100001110;
            15'd18835: log10_cal = 16'b0000010100001111;
            15'd18836: log10_cal = 16'b0000010100001111;
            15'd18837: log10_cal = 16'b0000010100001111;
            15'd18838: log10_cal = 16'b0000010100001111;
            15'd18839: log10_cal = 16'b0000010100001111;
            15'd18840: log10_cal = 16'b0000010100001111;
            15'd18841: log10_cal = 16'b0000010100001111;
            15'd18842: log10_cal = 16'b0000010100001111;
            15'd18843: log10_cal = 16'b0000010100001111;
            15'd18844: log10_cal = 16'b0000010100001111;
            15'd18845: log10_cal = 16'b0000010100001111;
            15'd18846: log10_cal = 16'b0000010100001111;
            15'd18847: log10_cal = 16'b0000010100001111;
            15'd18848: log10_cal = 16'b0000010100001111;
            15'd18849: log10_cal = 16'b0000010100001111;
            15'd18850: log10_cal = 16'b0000010100001111;
            15'd18851: log10_cal = 16'b0000010100001111;
            15'd18852: log10_cal = 16'b0000010100001111;
            15'd18853: log10_cal = 16'b0000010100001111;
            15'd18854: log10_cal = 16'b0000010100001111;
            15'd18855: log10_cal = 16'b0000010100001111;
            15'd18856: log10_cal = 16'b0000010100001111;
            15'd18857: log10_cal = 16'b0000010100001111;
            15'd18858: log10_cal = 16'b0000010100001111;
            15'd18859: log10_cal = 16'b0000010100001111;
            15'd18860: log10_cal = 16'b0000010100001111;
            15'd18861: log10_cal = 16'b0000010100001111;
            15'd18862: log10_cal = 16'b0000010100001111;
            15'd18863: log10_cal = 16'b0000010100001111;
            15'd18864: log10_cal = 16'b0000010100001111;
            15'd18865: log10_cal = 16'b0000010100001111;
            15'd18866: log10_cal = 16'b0000010100001111;
            15'd18867: log10_cal = 16'b0000010100001111;
            15'd18868: log10_cal = 16'b0000010100001111;
            15'd18869: log10_cal = 16'b0000010100001111;
            15'd18870: log10_cal = 16'b0000010100001111;
            15'd18871: log10_cal = 16'b0000010100001111;
            15'd18872: log10_cal = 16'b0000010100001111;
            15'd18873: log10_cal = 16'b0000010100001111;
            15'd18874: log10_cal = 16'b0000010100001111;
            15'd18875: log10_cal = 16'b0000010100001111;
            15'd18876: log10_cal = 16'b0000010100001111;
            15'd18877: log10_cal = 16'b0000010100010000;
            15'd18878: log10_cal = 16'b0000010100010000;
            15'd18879: log10_cal = 16'b0000010100010000;
            15'd18880: log10_cal = 16'b0000010100010000;
            15'd18881: log10_cal = 16'b0000010100010000;
            15'd18882: log10_cal = 16'b0000010100010000;
            15'd18883: log10_cal = 16'b0000010100010000;
            15'd18884: log10_cal = 16'b0000010100010000;
            15'd18885: log10_cal = 16'b0000010100010000;
            15'd18886: log10_cal = 16'b0000010100010000;
            15'd18887: log10_cal = 16'b0000010100010000;
            15'd18888: log10_cal = 16'b0000010100010000;
            15'd18889: log10_cal = 16'b0000010100010000;
            15'd18890: log10_cal = 16'b0000010100010000;
            15'd18891: log10_cal = 16'b0000010100010000;
            15'd18892: log10_cal = 16'b0000010100010000;
            15'd18893: log10_cal = 16'b0000010100010000;
            15'd18894: log10_cal = 16'b0000010100010000;
            15'd18895: log10_cal = 16'b0000010100010000;
            15'd18896: log10_cal = 16'b0000010100010000;
            15'd18897: log10_cal = 16'b0000010100010000;
            15'd18898: log10_cal = 16'b0000010100010000;
            15'd18899: log10_cal = 16'b0000010100010000;
            15'd18900: log10_cal = 16'b0000010100010000;
            15'd18901: log10_cal = 16'b0000010100010000;
            15'd18902: log10_cal = 16'b0000010100010000;
            15'd18903: log10_cal = 16'b0000010100010000;
            15'd18904: log10_cal = 16'b0000010100010000;
            15'd18905: log10_cal = 16'b0000010100010000;
            15'd18906: log10_cal = 16'b0000010100010000;
            15'd18907: log10_cal = 16'b0000010100010000;
            15'd18908: log10_cal = 16'b0000010100010000;
            15'd18909: log10_cal = 16'b0000010100010000;
            15'd18910: log10_cal = 16'b0000010100010000;
            15'd18911: log10_cal = 16'b0000010100010000;
            15'd18912: log10_cal = 16'b0000010100010000;
            15'd18913: log10_cal = 16'b0000010100010000;
            15'd18914: log10_cal = 16'b0000010100010000;
            15'd18915: log10_cal = 16'b0000010100010000;
            15'd18916: log10_cal = 16'b0000010100010000;
            15'd18917: log10_cal = 16'b0000010100010000;
            15'd18918: log10_cal = 16'b0000010100010000;
            15'd18919: log10_cal = 16'b0000010100010000;
            15'd18920: log10_cal = 16'b0000010100010001;
            15'd18921: log10_cal = 16'b0000010100010001;
            15'd18922: log10_cal = 16'b0000010100010001;
            15'd18923: log10_cal = 16'b0000010100010001;
            15'd18924: log10_cal = 16'b0000010100010001;
            15'd18925: log10_cal = 16'b0000010100010001;
            15'd18926: log10_cal = 16'b0000010100010001;
            15'd18927: log10_cal = 16'b0000010100010001;
            15'd18928: log10_cal = 16'b0000010100010001;
            15'd18929: log10_cal = 16'b0000010100010001;
            15'd18930: log10_cal = 16'b0000010100010001;
            15'd18931: log10_cal = 16'b0000010100010001;
            15'd18932: log10_cal = 16'b0000010100010001;
            15'd18933: log10_cal = 16'b0000010100010001;
            15'd18934: log10_cal = 16'b0000010100010001;
            15'd18935: log10_cal = 16'b0000010100010001;
            15'd18936: log10_cal = 16'b0000010100010001;
            15'd18937: log10_cal = 16'b0000010100010001;
            15'd18938: log10_cal = 16'b0000010100010001;
            15'd18939: log10_cal = 16'b0000010100010001;
            15'd18940: log10_cal = 16'b0000010100010001;
            15'd18941: log10_cal = 16'b0000010100010001;
            15'd18942: log10_cal = 16'b0000010100010001;
            15'd18943: log10_cal = 16'b0000010100010001;
            15'd18944: log10_cal = 16'b0000010100010001;
            15'd18945: log10_cal = 16'b0000010100010001;
            15'd18946: log10_cal = 16'b0000010100010001;
            15'd18947: log10_cal = 16'b0000010100010001;
            15'd18948: log10_cal = 16'b0000010100010001;
            15'd18949: log10_cal = 16'b0000010100010001;
            15'd18950: log10_cal = 16'b0000010100010001;
            15'd18951: log10_cal = 16'b0000010100010001;
            15'd18952: log10_cal = 16'b0000010100010001;
            15'd18953: log10_cal = 16'b0000010100010001;
            15'd18954: log10_cal = 16'b0000010100010001;
            15'd18955: log10_cal = 16'b0000010100010001;
            15'd18956: log10_cal = 16'b0000010100010001;
            15'd18957: log10_cal = 16'b0000010100010001;
            15'd18958: log10_cal = 16'b0000010100010001;
            15'd18959: log10_cal = 16'b0000010100010001;
            15'd18960: log10_cal = 16'b0000010100010001;
            15'd18961: log10_cal = 16'b0000010100010001;
            15'd18962: log10_cal = 16'b0000010100010010;
            15'd18963: log10_cal = 16'b0000010100010010;
            15'd18964: log10_cal = 16'b0000010100010010;
            15'd18965: log10_cal = 16'b0000010100010010;
            15'd18966: log10_cal = 16'b0000010100010010;
            15'd18967: log10_cal = 16'b0000010100010010;
            15'd18968: log10_cal = 16'b0000010100010010;
            15'd18969: log10_cal = 16'b0000010100010010;
            15'd18970: log10_cal = 16'b0000010100010010;
            15'd18971: log10_cal = 16'b0000010100010010;
            15'd18972: log10_cal = 16'b0000010100010010;
            15'd18973: log10_cal = 16'b0000010100010010;
            15'd18974: log10_cal = 16'b0000010100010010;
            15'd18975: log10_cal = 16'b0000010100010010;
            15'd18976: log10_cal = 16'b0000010100010010;
            15'd18977: log10_cal = 16'b0000010100010010;
            15'd18978: log10_cal = 16'b0000010100010010;
            15'd18979: log10_cal = 16'b0000010100010010;
            15'd18980: log10_cal = 16'b0000010100010010;
            15'd18981: log10_cal = 16'b0000010100010010;
            15'd18982: log10_cal = 16'b0000010100010010;
            15'd18983: log10_cal = 16'b0000010100010010;
            15'd18984: log10_cal = 16'b0000010100010010;
            15'd18985: log10_cal = 16'b0000010100010010;
            15'd18986: log10_cal = 16'b0000010100010010;
            15'd18987: log10_cal = 16'b0000010100010010;
            15'd18988: log10_cal = 16'b0000010100010010;
            15'd18989: log10_cal = 16'b0000010100010010;
            15'd18990: log10_cal = 16'b0000010100010010;
            15'd18991: log10_cal = 16'b0000010100010010;
            15'd18992: log10_cal = 16'b0000010100010010;
            15'd18993: log10_cal = 16'b0000010100010010;
            15'd18994: log10_cal = 16'b0000010100010010;
            15'd18995: log10_cal = 16'b0000010100010010;
            15'd18996: log10_cal = 16'b0000010100010010;
            15'd18997: log10_cal = 16'b0000010100010010;
            15'd18998: log10_cal = 16'b0000010100010010;
            15'd18999: log10_cal = 16'b0000010100010010;
            15'd19000: log10_cal = 16'b0000010100010010;
            15'd19001: log10_cal = 16'b0000010100010010;
            15'd19002: log10_cal = 16'b0000010100010010;
            15'd19003: log10_cal = 16'b0000010100010010;
            15'd19004: log10_cal = 16'b0000010100010010;
            15'd19005: log10_cal = 16'b0000010100010011;
            15'd19006: log10_cal = 16'b0000010100010011;
            15'd19007: log10_cal = 16'b0000010100010011;
            15'd19008: log10_cal = 16'b0000010100010011;
            15'd19009: log10_cal = 16'b0000010100010011;
            15'd19010: log10_cal = 16'b0000010100010011;
            15'd19011: log10_cal = 16'b0000010100010011;
            15'd19012: log10_cal = 16'b0000010100010011;
            15'd19013: log10_cal = 16'b0000010100010011;
            15'd19014: log10_cal = 16'b0000010100010011;
            15'd19015: log10_cal = 16'b0000010100010011;
            15'd19016: log10_cal = 16'b0000010100010011;
            15'd19017: log10_cal = 16'b0000010100010011;
            15'd19018: log10_cal = 16'b0000010100010011;
            15'd19019: log10_cal = 16'b0000010100010011;
            15'd19020: log10_cal = 16'b0000010100010011;
            15'd19021: log10_cal = 16'b0000010100010011;
            15'd19022: log10_cal = 16'b0000010100010011;
            15'd19023: log10_cal = 16'b0000010100010011;
            15'd19024: log10_cal = 16'b0000010100010011;
            15'd19025: log10_cal = 16'b0000010100010011;
            15'd19026: log10_cal = 16'b0000010100010011;
            15'd19027: log10_cal = 16'b0000010100010011;
            15'd19028: log10_cal = 16'b0000010100010011;
            15'd19029: log10_cal = 16'b0000010100010011;
            15'd19030: log10_cal = 16'b0000010100010011;
            15'd19031: log10_cal = 16'b0000010100010011;
            15'd19032: log10_cal = 16'b0000010100010011;
            15'd19033: log10_cal = 16'b0000010100010011;
            15'd19034: log10_cal = 16'b0000010100010011;
            15'd19035: log10_cal = 16'b0000010100010011;
            15'd19036: log10_cal = 16'b0000010100010011;
            15'd19037: log10_cal = 16'b0000010100010011;
            15'd19038: log10_cal = 16'b0000010100010011;
            15'd19039: log10_cal = 16'b0000010100010011;
            15'd19040: log10_cal = 16'b0000010100010011;
            15'd19041: log10_cal = 16'b0000010100010011;
            15'd19042: log10_cal = 16'b0000010100010011;
            15'd19043: log10_cal = 16'b0000010100010011;
            15'd19044: log10_cal = 16'b0000010100010011;
            15'd19045: log10_cal = 16'b0000010100010011;
            15'd19046: log10_cal = 16'b0000010100010011;
            15'd19047: log10_cal = 16'b0000010100010011;
            15'd19048: log10_cal = 16'b0000010100010100;
            15'd19049: log10_cal = 16'b0000010100010100;
            15'd19050: log10_cal = 16'b0000010100010100;
            15'd19051: log10_cal = 16'b0000010100010100;
            15'd19052: log10_cal = 16'b0000010100010100;
            15'd19053: log10_cal = 16'b0000010100010100;
            15'd19054: log10_cal = 16'b0000010100010100;
            15'd19055: log10_cal = 16'b0000010100010100;
            15'd19056: log10_cal = 16'b0000010100010100;
            15'd19057: log10_cal = 16'b0000010100010100;
            15'd19058: log10_cal = 16'b0000010100010100;
            15'd19059: log10_cal = 16'b0000010100010100;
            15'd19060: log10_cal = 16'b0000010100010100;
            15'd19061: log10_cal = 16'b0000010100010100;
            15'd19062: log10_cal = 16'b0000010100010100;
            15'd19063: log10_cal = 16'b0000010100010100;
            15'd19064: log10_cal = 16'b0000010100010100;
            15'd19065: log10_cal = 16'b0000010100010100;
            15'd19066: log10_cal = 16'b0000010100010100;
            15'd19067: log10_cal = 16'b0000010100010100;
            15'd19068: log10_cal = 16'b0000010100010100;
            15'd19069: log10_cal = 16'b0000010100010100;
            15'd19070: log10_cal = 16'b0000010100010100;
            15'd19071: log10_cal = 16'b0000010100010100;
            15'd19072: log10_cal = 16'b0000010100010100;
            15'd19073: log10_cal = 16'b0000010100010100;
            15'd19074: log10_cal = 16'b0000010100010100;
            15'd19075: log10_cal = 16'b0000010100010100;
            15'd19076: log10_cal = 16'b0000010100010100;
            15'd19077: log10_cal = 16'b0000010100010100;
            15'd19078: log10_cal = 16'b0000010100010100;
            15'd19079: log10_cal = 16'b0000010100010100;
            15'd19080: log10_cal = 16'b0000010100010100;
            15'd19081: log10_cal = 16'b0000010100010100;
            15'd19082: log10_cal = 16'b0000010100010100;
            15'd19083: log10_cal = 16'b0000010100010100;
            15'd19084: log10_cal = 16'b0000010100010100;
            15'd19085: log10_cal = 16'b0000010100010100;
            15'd19086: log10_cal = 16'b0000010100010100;
            15'd19087: log10_cal = 16'b0000010100010100;
            15'd19088: log10_cal = 16'b0000010100010100;
            15'd19089: log10_cal = 16'b0000010100010100;
            15'd19090: log10_cal = 16'b0000010100010100;
            15'd19091: log10_cal = 16'b0000010100010101;
            15'd19092: log10_cal = 16'b0000010100010101;
            15'd19093: log10_cal = 16'b0000010100010101;
            15'd19094: log10_cal = 16'b0000010100010101;
            15'd19095: log10_cal = 16'b0000010100010101;
            15'd19096: log10_cal = 16'b0000010100010101;
            15'd19097: log10_cal = 16'b0000010100010101;
            15'd19098: log10_cal = 16'b0000010100010101;
            15'd19099: log10_cal = 16'b0000010100010101;
            15'd19100: log10_cal = 16'b0000010100010101;
            15'd19101: log10_cal = 16'b0000010100010101;
            15'd19102: log10_cal = 16'b0000010100010101;
            15'd19103: log10_cal = 16'b0000010100010101;
            15'd19104: log10_cal = 16'b0000010100010101;
            15'd19105: log10_cal = 16'b0000010100010101;
            15'd19106: log10_cal = 16'b0000010100010101;
            15'd19107: log10_cal = 16'b0000010100010101;
            15'd19108: log10_cal = 16'b0000010100010101;
            15'd19109: log10_cal = 16'b0000010100010101;
            15'd19110: log10_cal = 16'b0000010100010101;
            15'd19111: log10_cal = 16'b0000010100010101;
            15'd19112: log10_cal = 16'b0000010100010101;
            15'd19113: log10_cal = 16'b0000010100010101;
            15'd19114: log10_cal = 16'b0000010100010101;
            15'd19115: log10_cal = 16'b0000010100010101;
            15'd19116: log10_cal = 16'b0000010100010101;
            15'd19117: log10_cal = 16'b0000010100010101;
            15'd19118: log10_cal = 16'b0000010100010101;
            15'd19119: log10_cal = 16'b0000010100010101;
            15'd19120: log10_cal = 16'b0000010100010101;
            15'd19121: log10_cal = 16'b0000010100010101;
            15'd19122: log10_cal = 16'b0000010100010101;
            15'd19123: log10_cal = 16'b0000010100010101;
            15'd19124: log10_cal = 16'b0000010100010101;
            15'd19125: log10_cal = 16'b0000010100010101;
            15'd19126: log10_cal = 16'b0000010100010101;
            15'd19127: log10_cal = 16'b0000010100010101;
            15'd19128: log10_cal = 16'b0000010100010101;
            15'd19129: log10_cal = 16'b0000010100010101;
            15'd19130: log10_cal = 16'b0000010100010101;
            15'd19131: log10_cal = 16'b0000010100010101;
            15'd19132: log10_cal = 16'b0000010100010101;
            15'd19133: log10_cal = 16'b0000010100010101;
            15'd19134: log10_cal = 16'b0000010100010110;
            15'd19135: log10_cal = 16'b0000010100010110;
            15'd19136: log10_cal = 16'b0000010100010110;
            15'd19137: log10_cal = 16'b0000010100010110;
            15'd19138: log10_cal = 16'b0000010100010110;
            15'd19139: log10_cal = 16'b0000010100010110;
            15'd19140: log10_cal = 16'b0000010100010110;
            15'd19141: log10_cal = 16'b0000010100010110;
            15'd19142: log10_cal = 16'b0000010100010110;
            15'd19143: log10_cal = 16'b0000010100010110;
            15'd19144: log10_cal = 16'b0000010100010110;
            15'd19145: log10_cal = 16'b0000010100010110;
            15'd19146: log10_cal = 16'b0000010100010110;
            15'd19147: log10_cal = 16'b0000010100010110;
            15'd19148: log10_cal = 16'b0000010100010110;
            15'd19149: log10_cal = 16'b0000010100010110;
            15'd19150: log10_cal = 16'b0000010100010110;
            15'd19151: log10_cal = 16'b0000010100010110;
            15'd19152: log10_cal = 16'b0000010100010110;
            15'd19153: log10_cal = 16'b0000010100010110;
            15'd19154: log10_cal = 16'b0000010100010110;
            15'd19155: log10_cal = 16'b0000010100010110;
            15'd19156: log10_cal = 16'b0000010100010110;
            15'd19157: log10_cal = 16'b0000010100010110;
            15'd19158: log10_cal = 16'b0000010100010110;
            15'd19159: log10_cal = 16'b0000010100010110;
            15'd19160: log10_cal = 16'b0000010100010110;
            15'd19161: log10_cal = 16'b0000010100010110;
            15'd19162: log10_cal = 16'b0000010100010110;
            15'd19163: log10_cal = 16'b0000010100010110;
            15'd19164: log10_cal = 16'b0000010100010110;
            15'd19165: log10_cal = 16'b0000010100010110;
            15'd19166: log10_cal = 16'b0000010100010110;
            15'd19167: log10_cal = 16'b0000010100010110;
            15'd19168: log10_cal = 16'b0000010100010110;
            15'd19169: log10_cal = 16'b0000010100010110;
            15'd19170: log10_cal = 16'b0000010100010110;
            15'd19171: log10_cal = 16'b0000010100010110;
            15'd19172: log10_cal = 16'b0000010100010110;
            15'd19173: log10_cal = 16'b0000010100010110;
            15'd19174: log10_cal = 16'b0000010100010110;
            15'd19175: log10_cal = 16'b0000010100010110;
            15'd19176: log10_cal = 16'b0000010100010110;
            15'd19177: log10_cal = 16'b0000010100010111;
            15'd19178: log10_cal = 16'b0000010100010111;
            15'd19179: log10_cal = 16'b0000010100010111;
            15'd19180: log10_cal = 16'b0000010100010111;
            15'd19181: log10_cal = 16'b0000010100010111;
            15'd19182: log10_cal = 16'b0000010100010111;
            15'd19183: log10_cal = 16'b0000010100010111;
            15'd19184: log10_cal = 16'b0000010100010111;
            15'd19185: log10_cal = 16'b0000010100010111;
            15'd19186: log10_cal = 16'b0000010100010111;
            15'd19187: log10_cal = 16'b0000010100010111;
            15'd19188: log10_cal = 16'b0000010100010111;
            15'd19189: log10_cal = 16'b0000010100010111;
            15'd19190: log10_cal = 16'b0000010100010111;
            15'd19191: log10_cal = 16'b0000010100010111;
            15'd19192: log10_cal = 16'b0000010100010111;
            15'd19193: log10_cal = 16'b0000010100010111;
            15'd19194: log10_cal = 16'b0000010100010111;
            15'd19195: log10_cal = 16'b0000010100010111;
            15'd19196: log10_cal = 16'b0000010100010111;
            15'd19197: log10_cal = 16'b0000010100010111;
            15'd19198: log10_cal = 16'b0000010100010111;
            15'd19199: log10_cal = 16'b0000010100010111;
            15'd19200: log10_cal = 16'b0000010100010111;
            15'd19201: log10_cal = 16'b0000010100010111;
            15'd19202: log10_cal = 16'b0000010100010111;
            15'd19203: log10_cal = 16'b0000010100010111;
            15'd19204: log10_cal = 16'b0000010100010111;
            15'd19205: log10_cal = 16'b0000010100010111;
            15'd19206: log10_cal = 16'b0000010100010111;
            15'd19207: log10_cal = 16'b0000010100010111;
            15'd19208: log10_cal = 16'b0000010100010111;
            15'd19209: log10_cal = 16'b0000010100010111;
            15'd19210: log10_cal = 16'b0000010100010111;
            15'd19211: log10_cal = 16'b0000010100010111;
            15'd19212: log10_cal = 16'b0000010100010111;
            15'd19213: log10_cal = 16'b0000010100010111;
            15'd19214: log10_cal = 16'b0000010100010111;
            15'd19215: log10_cal = 16'b0000010100010111;
            15'd19216: log10_cal = 16'b0000010100010111;
            15'd19217: log10_cal = 16'b0000010100010111;
            15'd19218: log10_cal = 16'b0000010100010111;
            15'd19219: log10_cal = 16'b0000010100010111;
            15'd19220: log10_cal = 16'b0000010100011000;
            15'd19221: log10_cal = 16'b0000010100011000;
            15'd19222: log10_cal = 16'b0000010100011000;
            15'd19223: log10_cal = 16'b0000010100011000;
            15'd19224: log10_cal = 16'b0000010100011000;
            15'd19225: log10_cal = 16'b0000010100011000;
            15'd19226: log10_cal = 16'b0000010100011000;
            15'd19227: log10_cal = 16'b0000010100011000;
            15'd19228: log10_cal = 16'b0000010100011000;
            15'd19229: log10_cal = 16'b0000010100011000;
            15'd19230: log10_cal = 16'b0000010100011000;
            15'd19231: log10_cal = 16'b0000010100011000;
            15'd19232: log10_cal = 16'b0000010100011000;
            15'd19233: log10_cal = 16'b0000010100011000;
            15'd19234: log10_cal = 16'b0000010100011000;
            15'd19235: log10_cal = 16'b0000010100011000;
            15'd19236: log10_cal = 16'b0000010100011000;
            15'd19237: log10_cal = 16'b0000010100011000;
            15'd19238: log10_cal = 16'b0000010100011000;
            15'd19239: log10_cal = 16'b0000010100011000;
            15'd19240: log10_cal = 16'b0000010100011000;
            15'd19241: log10_cal = 16'b0000010100011000;
            15'd19242: log10_cal = 16'b0000010100011000;
            15'd19243: log10_cal = 16'b0000010100011000;
            15'd19244: log10_cal = 16'b0000010100011000;
            15'd19245: log10_cal = 16'b0000010100011000;
            15'd19246: log10_cal = 16'b0000010100011000;
            15'd19247: log10_cal = 16'b0000010100011000;
            15'd19248: log10_cal = 16'b0000010100011000;
            15'd19249: log10_cal = 16'b0000010100011000;
            15'd19250: log10_cal = 16'b0000010100011000;
            15'd19251: log10_cal = 16'b0000010100011000;
            15'd19252: log10_cal = 16'b0000010100011000;
            15'd19253: log10_cal = 16'b0000010100011000;
            15'd19254: log10_cal = 16'b0000010100011000;
            15'd19255: log10_cal = 16'b0000010100011000;
            15'd19256: log10_cal = 16'b0000010100011000;
            15'd19257: log10_cal = 16'b0000010100011000;
            15'd19258: log10_cal = 16'b0000010100011000;
            15'd19259: log10_cal = 16'b0000010100011000;
            15'd19260: log10_cal = 16'b0000010100011000;
            15'd19261: log10_cal = 16'b0000010100011000;
            15'd19262: log10_cal = 16'b0000010100011000;
            15'd19263: log10_cal = 16'b0000010100011001;
            15'd19264: log10_cal = 16'b0000010100011001;
            15'd19265: log10_cal = 16'b0000010100011001;
            15'd19266: log10_cal = 16'b0000010100011001;
            15'd19267: log10_cal = 16'b0000010100011001;
            15'd19268: log10_cal = 16'b0000010100011001;
            15'd19269: log10_cal = 16'b0000010100011001;
            15'd19270: log10_cal = 16'b0000010100011001;
            15'd19271: log10_cal = 16'b0000010100011001;
            15'd19272: log10_cal = 16'b0000010100011001;
            15'd19273: log10_cal = 16'b0000010100011001;
            15'd19274: log10_cal = 16'b0000010100011001;
            15'd19275: log10_cal = 16'b0000010100011001;
            15'd19276: log10_cal = 16'b0000010100011001;
            15'd19277: log10_cal = 16'b0000010100011001;
            15'd19278: log10_cal = 16'b0000010100011001;
            15'd19279: log10_cal = 16'b0000010100011001;
            15'd19280: log10_cal = 16'b0000010100011001;
            15'd19281: log10_cal = 16'b0000010100011001;
            15'd19282: log10_cal = 16'b0000010100011001;
            15'd19283: log10_cal = 16'b0000010100011001;
            15'd19284: log10_cal = 16'b0000010100011001;
            15'd19285: log10_cal = 16'b0000010100011001;
            15'd19286: log10_cal = 16'b0000010100011001;
            15'd19287: log10_cal = 16'b0000010100011001;
            15'd19288: log10_cal = 16'b0000010100011001;
            15'd19289: log10_cal = 16'b0000010100011001;
            15'd19290: log10_cal = 16'b0000010100011001;
            15'd19291: log10_cal = 16'b0000010100011001;
            15'd19292: log10_cal = 16'b0000010100011001;
            15'd19293: log10_cal = 16'b0000010100011001;
            15'd19294: log10_cal = 16'b0000010100011001;
            15'd19295: log10_cal = 16'b0000010100011001;
            15'd19296: log10_cal = 16'b0000010100011001;
            15'd19297: log10_cal = 16'b0000010100011001;
            15'd19298: log10_cal = 16'b0000010100011001;
            15'd19299: log10_cal = 16'b0000010100011001;
            15'd19300: log10_cal = 16'b0000010100011001;
            15'd19301: log10_cal = 16'b0000010100011001;
            15'd19302: log10_cal = 16'b0000010100011001;
            15'd19303: log10_cal = 16'b0000010100011001;
            15'd19304: log10_cal = 16'b0000010100011001;
            15'd19305: log10_cal = 16'b0000010100011001;
            15'd19306: log10_cal = 16'b0000010100011010;
            15'd19307: log10_cal = 16'b0000010100011010;
            15'd19308: log10_cal = 16'b0000010100011010;
            15'd19309: log10_cal = 16'b0000010100011010;
            15'd19310: log10_cal = 16'b0000010100011010;
            15'd19311: log10_cal = 16'b0000010100011010;
            15'd19312: log10_cal = 16'b0000010100011010;
            15'd19313: log10_cal = 16'b0000010100011010;
            15'd19314: log10_cal = 16'b0000010100011010;
            15'd19315: log10_cal = 16'b0000010100011010;
            15'd19316: log10_cal = 16'b0000010100011010;
            15'd19317: log10_cal = 16'b0000010100011010;
            15'd19318: log10_cal = 16'b0000010100011010;
            15'd19319: log10_cal = 16'b0000010100011010;
            15'd19320: log10_cal = 16'b0000010100011010;
            15'd19321: log10_cal = 16'b0000010100011010;
            15'd19322: log10_cal = 16'b0000010100011010;
            15'd19323: log10_cal = 16'b0000010100011010;
            15'd19324: log10_cal = 16'b0000010100011010;
            15'd19325: log10_cal = 16'b0000010100011010;
            15'd19326: log10_cal = 16'b0000010100011010;
            15'd19327: log10_cal = 16'b0000010100011010;
            15'd19328: log10_cal = 16'b0000010100011010;
            15'd19329: log10_cal = 16'b0000010100011010;
            15'd19330: log10_cal = 16'b0000010100011010;
            15'd19331: log10_cal = 16'b0000010100011010;
            15'd19332: log10_cal = 16'b0000010100011010;
            15'd19333: log10_cal = 16'b0000010100011010;
            15'd19334: log10_cal = 16'b0000010100011010;
            15'd19335: log10_cal = 16'b0000010100011010;
            15'd19336: log10_cal = 16'b0000010100011010;
            15'd19337: log10_cal = 16'b0000010100011010;
            15'd19338: log10_cal = 16'b0000010100011010;
            15'd19339: log10_cal = 16'b0000010100011010;
            15'd19340: log10_cal = 16'b0000010100011010;
            15'd19341: log10_cal = 16'b0000010100011010;
            15'd19342: log10_cal = 16'b0000010100011010;
            15'd19343: log10_cal = 16'b0000010100011010;
            15'd19344: log10_cal = 16'b0000010100011010;
            15'd19345: log10_cal = 16'b0000010100011010;
            15'd19346: log10_cal = 16'b0000010100011010;
            15'd19347: log10_cal = 16'b0000010100011010;
            15'd19348: log10_cal = 16'b0000010100011010;
            15'd19349: log10_cal = 16'b0000010100011010;
            15'd19350: log10_cal = 16'b0000010100011011;
            15'd19351: log10_cal = 16'b0000010100011011;
            15'd19352: log10_cal = 16'b0000010100011011;
            15'd19353: log10_cal = 16'b0000010100011011;
            15'd19354: log10_cal = 16'b0000010100011011;
            15'd19355: log10_cal = 16'b0000010100011011;
            15'd19356: log10_cal = 16'b0000010100011011;
            15'd19357: log10_cal = 16'b0000010100011011;
            15'd19358: log10_cal = 16'b0000010100011011;
            15'd19359: log10_cal = 16'b0000010100011011;
            15'd19360: log10_cal = 16'b0000010100011011;
            15'd19361: log10_cal = 16'b0000010100011011;
            15'd19362: log10_cal = 16'b0000010100011011;
            15'd19363: log10_cal = 16'b0000010100011011;
            15'd19364: log10_cal = 16'b0000010100011011;
            15'd19365: log10_cal = 16'b0000010100011011;
            15'd19366: log10_cal = 16'b0000010100011011;
            15'd19367: log10_cal = 16'b0000010100011011;
            15'd19368: log10_cal = 16'b0000010100011011;
            15'd19369: log10_cal = 16'b0000010100011011;
            15'd19370: log10_cal = 16'b0000010100011011;
            15'd19371: log10_cal = 16'b0000010100011011;
            15'd19372: log10_cal = 16'b0000010100011011;
            15'd19373: log10_cal = 16'b0000010100011011;
            15'd19374: log10_cal = 16'b0000010100011011;
            15'd19375: log10_cal = 16'b0000010100011011;
            15'd19376: log10_cal = 16'b0000010100011011;
            15'd19377: log10_cal = 16'b0000010100011011;
            15'd19378: log10_cal = 16'b0000010100011011;
            15'd19379: log10_cal = 16'b0000010100011011;
            15'd19380: log10_cal = 16'b0000010100011011;
            15'd19381: log10_cal = 16'b0000010100011011;
            15'd19382: log10_cal = 16'b0000010100011011;
            15'd19383: log10_cal = 16'b0000010100011011;
            15'd19384: log10_cal = 16'b0000010100011011;
            15'd19385: log10_cal = 16'b0000010100011011;
            15'd19386: log10_cal = 16'b0000010100011011;
            15'd19387: log10_cal = 16'b0000010100011011;
            15'd19388: log10_cal = 16'b0000010100011011;
            15'd19389: log10_cal = 16'b0000010100011011;
            15'd19390: log10_cal = 16'b0000010100011011;
            15'd19391: log10_cal = 16'b0000010100011011;
            15'd19392: log10_cal = 16'b0000010100011011;
            15'd19393: log10_cal = 16'b0000010100011100;
            15'd19394: log10_cal = 16'b0000010100011100;
            15'd19395: log10_cal = 16'b0000010100011100;
            15'd19396: log10_cal = 16'b0000010100011100;
            15'd19397: log10_cal = 16'b0000010100011100;
            15'd19398: log10_cal = 16'b0000010100011100;
            15'd19399: log10_cal = 16'b0000010100011100;
            15'd19400: log10_cal = 16'b0000010100011100;
            15'd19401: log10_cal = 16'b0000010100011100;
            15'd19402: log10_cal = 16'b0000010100011100;
            15'd19403: log10_cal = 16'b0000010100011100;
            15'd19404: log10_cal = 16'b0000010100011100;
            15'd19405: log10_cal = 16'b0000010100011100;
            15'd19406: log10_cal = 16'b0000010100011100;
            15'd19407: log10_cal = 16'b0000010100011100;
            15'd19408: log10_cal = 16'b0000010100011100;
            15'd19409: log10_cal = 16'b0000010100011100;
            15'd19410: log10_cal = 16'b0000010100011100;
            15'd19411: log10_cal = 16'b0000010100011100;
            15'd19412: log10_cal = 16'b0000010100011100;
            15'd19413: log10_cal = 16'b0000010100011100;
            15'd19414: log10_cal = 16'b0000010100011100;
            15'd19415: log10_cal = 16'b0000010100011100;
            15'd19416: log10_cal = 16'b0000010100011100;
            15'd19417: log10_cal = 16'b0000010100011100;
            15'd19418: log10_cal = 16'b0000010100011100;
            15'd19419: log10_cal = 16'b0000010100011100;
            15'd19420: log10_cal = 16'b0000010100011100;
            15'd19421: log10_cal = 16'b0000010100011100;
            15'd19422: log10_cal = 16'b0000010100011100;
            15'd19423: log10_cal = 16'b0000010100011100;
            15'd19424: log10_cal = 16'b0000010100011100;
            15'd19425: log10_cal = 16'b0000010100011100;
            15'd19426: log10_cal = 16'b0000010100011100;
            15'd19427: log10_cal = 16'b0000010100011100;
            15'd19428: log10_cal = 16'b0000010100011100;
            15'd19429: log10_cal = 16'b0000010100011100;
            15'd19430: log10_cal = 16'b0000010100011100;
            15'd19431: log10_cal = 16'b0000010100011100;
            15'd19432: log10_cal = 16'b0000010100011100;
            15'd19433: log10_cal = 16'b0000010100011100;
            15'd19434: log10_cal = 16'b0000010100011100;
            15'd19435: log10_cal = 16'b0000010100011100;
            15'd19436: log10_cal = 16'b0000010100011100;
            15'd19437: log10_cal = 16'b0000010100011101;
            15'd19438: log10_cal = 16'b0000010100011101;
            15'd19439: log10_cal = 16'b0000010100011101;
            15'd19440: log10_cal = 16'b0000010100011101;
            15'd19441: log10_cal = 16'b0000010100011101;
            15'd19442: log10_cal = 16'b0000010100011101;
            15'd19443: log10_cal = 16'b0000010100011101;
            15'd19444: log10_cal = 16'b0000010100011101;
            15'd19445: log10_cal = 16'b0000010100011101;
            15'd19446: log10_cal = 16'b0000010100011101;
            15'd19447: log10_cal = 16'b0000010100011101;
            15'd19448: log10_cal = 16'b0000010100011101;
            15'd19449: log10_cal = 16'b0000010100011101;
            15'd19450: log10_cal = 16'b0000010100011101;
            15'd19451: log10_cal = 16'b0000010100011101;
            15'd19452: log10_cal = 16'b0000010100011101;
            15'd19453: log10_cal = 16'b0000010100011101;
            15'd19454: log10_cal = 16'b0000010100011101;
            15'd19455: log10_cal = 16'b0000010100011101;
            15'd19456: log10_cal = 16'b0000010100011101;
            15'd19457: log10_cal = 16'b0000010100011101;
            15'd19458: log10_cal = 16'b0000010100011101;
            15'd19459: log10_cal = 16'b0000010100011101;
            15'd19460: log10_cal = 16'b0000010100011101;
            15'd19461: log10_cal = 16'b0000010100011101;
            15'd19462: log10_cal = 16'b0000010100011101;
            15'd19463: log10_cal = 16'b0000010100011101;
            15'd19464: log10_cal = 16'b0000010100011101;
            15'd19465: log10_cal = 16'b0000010100011101;
            15'd19466: log10_cal = 16'b0000010100011101;
            15'd19467: log10_cal = 16'b0000010100011101;
            15'd19468: log10_cal = 16'b0000010100011101;
            15'd19469: log10_cal = 16'b0000010100011101;
            15'd19470: log10_cal = 16'b0000010100011101;
            15'd19471: log10_cal = 16'b0000010100011101;
            15'd19472: log10_cal = 16'b0000010100011101;
            15'd19473: log10_cal = 16'b0000010100011101;
            15'd19474: log10_cal = 16'b0000010100011101;
            15'd19475: log10_cal = 16'b0000010100011101;
            15'd19476: log10_cal = 16'b0000010100011101;
            15'd19477: log10_cal = 16'b0000010100011101;
            15'd19478: log10_cal = 16'b0000010100011101;
            15'd19479: log10_cal = 16'b0000010100011101;
            15'd19480: log10_cal = 16'b0000010100011101;
            15'd19481: log10_cal = 16'b0000010100011110;
            15'd19482: log10_cal = 16'b0000010100011110;
            15'd19483: log10_cal = 16'b0000010100011110;
            15'd19484: log10_cal = 16'b0000010100011110;
            15'd19485: log10_cal = 16'b0000010100011110;
            15'd19486: log10_cal = 16'b0000010100011110;
            15'd19487: log10_cal = 16'b0000010100011110;
            15'd19488: log10_cal = 16'b0000010100011110;
            15'd19489: log10_cal = 16'b0000010100011110;
            15'd19490: log10_cal = 16'b0000010100011110;
            15'd19491: log10_cal = 16'b0000010100011110;
            15'd19492: log10_cal = 16'b0000010100011110;
            15'd19493: log10_cal = 16'b0000010100011110;
            15'd19494: log10_cal = 16'b0000010100011110;
            15'd19495: log10_cal = 16'b0000010100011110;
            15'd19496: log10_cal = 16'b0000010100011110;
            15'd19497: log10_cal = 16'b0000010100011110;
            15'd19498: log10_cal = 16'b0000010100011110;
            15'd19499: log10_cal = 16'b0000010100011110;
            15'd19500: log10_cal = 16'b0000010100011110;
            15'd19501: log10_cal = 16'b0000010100011110;
            15'd19502: log10_cal = 16'b0000010100011110;
            15'd19503: log10_cal = 16'b0000010100011110;
            15'd19504: log10_cal = 16'b0000010100011110;
            15'd19505: log10_cal = 16'b0000010100011110;
            15'd19506: log10_cal = 16'b0000010100011110;
            15'd19507: log10_cal = 16'b0000010100011110;
            15'd19508: log10_cal = 16'b0000010100011110;
            15'd19509: log10_cal = 16'b0000010100011110;
            15'd19510: log10_cal = 16'b0000010100011110;
            15'd19511: log10_cal = 16'b0000010100011110;
            15'd19512: log10_cal = 16'b0000010100011110;
            15'd19513: log10_cal = 16'b0000010100011110;
            15'd19514: log10_cal = 16'b0000010100011110;
            15'd19515: log10_cal = 16'b0000010100011110;
            15'd19516: log10_cal = 16'b0000010100011110;
            15'd19517: log10_cal = 16'b0000010100011110;
            15'd19518: log10_cal = 16'b0000010100011110;
            15'd19519: log10_cal = 16'b0000010100011110;
            15'd19520: log10_cal = 16'b0000010100011110;
            15'd19521: log10_cal = 16'b0000010100011110;
            15'd19522: log10_cal = 16'b0000010100011110;
            15'd19523: log10_cal = 16'b0000010100011110;
            15'd19524: log10_cal = 16'b0000010100011110;
            15'd19525: log10_cal = 16'b0000010100011111;
            15'd19526: log10_cal = 16'b0000010100011111;
            15'd19527: log10_cal = 16'b0000010100011111;
            15'd19528: log10_cal = 16'b0000010100011111;
            15'd19529: log10_cal = 16'b0000010100011111;
            15'd19530: log10_cal = 16'b0000010100011111;
            15'd19531: log10_cal = 16'b0000010100011111;
            15'd19532: log10_cal = 16'b0000010100011111;
            15'd19533: log10_cal = 16'b0000010100011111;
            15'd19534: log10_cal = 16'b0000010100011111;
            15'd19535: log10_cal = 16'b0000010100011111;
            15'd19536: log10_cal = 16'b0000010100011111;
            15'd19537: log10_cal = 16'b0000010100011111;
            15'd19538: log10_cal = 16'b0000010100011111;
            15'd19539: log10_cal = 16'b0000010100011111;
            15'd19540: log10_cal = 16'b0000010100011111;
            15'd19541: log10_cal = 16'b0000010100011111;
            15'd19542: log10_cal = 16'b0000010100011111;
            15'd19543: log10_cal = 16'b0000010100011111;
            15'd19544: log10_cal = 16'b0000010100011111;
            15'd19545: log10_cal = 16'b0000010100011111;
            15'd19546: log10_cal = 16'b0000010100011111;
            15'd19547: log10_cal = 16'b0000010100011111;
            15'd19548: log10_cal = 16'b0000010100011111;
            15'd19549: log10_cal = 16'b0000010100011111;
            15'd19550: log10_cal = 16'b0000010100011111;
            15'd19551: log10_cal = 16'b0000010100011111;
            15'd19552: log10_cal = 16'b0000010100011111;
            15'd19553: log10_cal = 16'b0000010100011111;
            15'd19554: log10_cal = 16'b0000010100011111;
            15'd19555: log10_cal = 16'b0000010100011111;
            15'd19556: log10_cal = 16'b0000010100011111;
            15'd19557: log10_cal = 16'b0000010100011111;
            15'd19558: log10_cal = 16'b0000010100011111;
            15'd19559: log10_cal = 16'b0000010100011111;
            15'd19560: log10_cal = 16'b0000010100011111;
            15'd19561: log10_cal = 16'b0000010100011111;
            15'd19562: log10_cal = 16'b0000010100011111;
            15'd19563: log10_cal = 16'b0000010100011111;
            15'd19564: log10_cal = 16'b0000010100011111;
            15'd19565: log10_cal = 16'b0000010100011111;
            15'd19566: log10_cal = 16'b0000010100011111;
            15'd19567: log10_cal = 16'b0000010100011111;
            15'd19568: log10_cal = 16'b0000010100011111;
            15'd19569: log10_cal = 16'b0000010100100000;
            15'd19570: log10_cal = 16'b0000010100100000;
            15'd19571: log10_cal = 16'b0000010100100000;
            15'd19572: log10_cal = 16'b0000010100100000;
            15'd19573: log10_cal = 16'b0000010100100000;
            15'd19574: log10_cal = 16'b0000010100100000;
            15'd19575: log10_cal = 16'b0000010100100000;
            15'd19576: log10_cal = 16'b0000010100100000;
            15'd19577: log10_cal = 16'b0000010100100000;
            15'd19578: log10_cal = 16'b0000010100100000;
            15'd19579: log10_cal = 16'b0000010100100000;
            15'd19580: log10_cal = 16'b0000010100100000;
            15'd19581: log10_cal = 16'b0000010100100000;
            15'd19582: log10_cal = 16'b0000010100100000;
            15'd19583: log10_cal = 16'b0000010100100000;
            15'd19584: log10_cal = 16'b0000010100100000;
            15'd19585: log10_cal = 16'b0000010100100000;
            15'd19586: log10_cal = 16'b0000010100100000;
            15'd19587: log10_cal = 16'b0000010100100000;
            15'd19588: log10_cal = 16'b0000010100100000;
            15'd19589: log10_cal = 16'b0000010100100000;
            15'd19590: log10_cal = 16'b0000010100100000;
            15'd19591: log10_cal = 16'b0000010100100000;
            15'd19592: log10_cal = 16'b0000010100100000;
            15'd19593: log10_cal = 16'b0000010100100000;
            15'd19594: log10_cal = 16'b0000010100100000;
            15'd19595: log10_cal = 16'b0000010100100000;
            15'd19596: log10_cal = 16'b0000010100100000;
            15'd19597: log10_cal = 16'b0000010100100000;
            15'd19598: log10_cal = 16'b0000010100100000;
            15'd19599: log10_cal = 16'b0000010100100000;
            15'd19600: log10_cal = 16'b0000010100100000;
            15'd19601: log10_cal = 16'b0000010100100000;
            15'd19602: log10_cal = 16'b0000010100100000;
            15'd19603: log10_cal = 16'b0000010100100000;
            15'd19604: log10_cal = 16'b0000010100100000;
            15'd19605: log10_cal = 16'b0000010100100000;
            15'd19606: log10_cal = 16'b0000010100100000;
            15'd19607: log10_cal = 16'b0000010100100000;
            15'd19608: log10_cal = 16'b0000010100100000;
            15'd19609: log10_cal = 16'b0000010100100000;
            15'd19610: log10_cal = 16'b0000010100100000;
            15'd19611: log10_cal = 16'b0000010100100000;
            15'd19612: log10_cal = 16'b0000010100100000;
            15'd19613: log10_cal = 16'b0000010100100001;
            15'd19614: log10_cal = 16'b0000010100100001;
            15'd19615: log10_cal = 16'b0000010100100001;
            15'd19616: log10_cal = 16'b0000010100100001;
            15'd19617: log10_cal = 16'b0000010100100001;
            15'd19618: log10_cal = 16'b0000010100100001;
            15'd19619: log10_cal = 16'b0000010100100001;
            15'd19620: log10_cal = 16'b0000010100100001;
            15'd19621: log10_cal = 16'b0000010100100001;
            15'd19622: log10_cal = 16'b0000010100100001;
            15'd19623: log10_cal = 16'b0000010100100001;
            15'd19624: log10_cal = 16'b0000010100100001;
            15'd19625: log10_cal = 16'b0000010100100001;
            15'd19626: log10_cal = 16'b0000010100100001;
            15'd19627: log10_cal = 16'b0000010100100001;
            15'd19628: log10_cal = 16'b0000010100100001;
            15'd19629: log10_cal = 16'b0000010100100001;
            15'd19630: log10_cal = 16'b0000010100100001;
            15'd19631: log10_cal = 16'b0000010100100001;
            15'd19632: log10_cal = 16'b0000010100100001;
            15'd19633: log10_cal = 16'b0000010100100001;
            15'd19634: log10_cal = 16'b0000010100100001;
            15'd19635: log10_cal = 16'b0000010100100001;
            15'd19636: log10_cal = 16'b0000010100100001;
            15'd19637: log10_cal = 16'b0000010100100001;
            15'd19638: log10_cal = 16'b0000010100100001;
            15'd19639: log10_cal = 16'b0000010100100001;
            15'd19640: log10_cal = 16'b0000010100100001;
            15'd19641: log10_cal = 16'b0000010100100001;
            15'd19642: log10_cal = 16'b0000010100100001;
            15'd19643: log10_cal = 16'b0000010100100001;
            15'd19644: log10_cal = 16'b0000010100100001;
            15'd19645: log10_cal = 16'b0000010100100001;
            15'd19646: log10_cal = 16'b0000010100100001;
            15'd19647: log10_cal = 16'b0000010100100001;
            15'd19648: log10_cal = 16'b0000010100100001;
            15'd19649: log10_cal = 16'b0000010100100001;
            15'd19650: log10_cal = 16'b0000010100100001;
            15'd19651: log10_cal = 16'b0000010100100001;
            15'd19652: log10_cal = 16'b0000010100100001;
            15'd19653: log10_cal = 16'b0000010100100001;
            15'd19654: log10_cal = 16'b0000010100100001;
            15'd19655: log10_cal = 16'b0000010100100001;
            15'd19656: log10_cal = 16'b0000010100100001;
            15'd19657: log10_cal = 16'b0000010100100010;
            15'd19658: log10_cal = 16'b0000010100100010;
            15'd19659: log10_cal = 16'b0000010100100010;
            15'd19660: log10_cal = 16'b0000010100100010;
            15'd19661: log10_cal = 16'b0000010100100010;
            15'd19662: log10_cal = 16'b0000010100100010;
            15'd19663: log10_cal = 16'b0000010100100010;
            15'd19664: log10_cal = 16'b0000010100100010;
            15'd19665: log10_cal = 16'b0000010100100010;
            15'd19666: log10_cal = 16'b0000010100100010;
            15'd19667: log10_cal = 16'b0000010100100010;
            15'd19668: log10_cal = 16'b0000010100100010;
            15'd19669: log10_cal = 16'b0000010100100010;
            15'd19670: log10_cal = 16'b0000010100100010;
            15'd19671: log10_cal = 16'b0000010100100010;
            15'd19672: log10_cal = 16'b0000010100100010;
            15'd19673: log10_cal = 16'b0000010100100010;
            15'd19674: log10_cal = 16'b0000010100100010;
            15'd19675: log10_cal = 16'b0000010100100010;
            15'd19676: log10_cal = 16'b0000010100100010;
            15'd19677: log10_cal = 16'b0000010100100010;
            15'd19678: log10_cal = 16'b0000010100100010;
            15'd19679: log10_cal = 16'b0000010100100010;
            15'd19680: log10_cal = 16'b0000010100100010;
            15'd19681: log10_cal = 16'b0000010100100010;
            15'd19682: log10_cal = 16'b0000010100100010;
            15'd19683: log10_cal = 16'b0000010100100010;
            15'd19684: log10_cal = 16'b0000010100100010;
            15'd19685: log10_cal = 16'b0000010100100010;
            15'd19686: log10_cal = 16'b0000010100100010;
            15'd19687: log10_cal = 16'b0000010100100010;
            15'd19688: log10_cal = 16'b0000010100100010;
            15'd19689: log10_cal = 16'b0000010100100010;
            15'd19690: log10_cal = 16'b0000010100100010;
            15'd19691: log10_cal = 16'b0000010100100010;
            15'd19692: log10_cal = 16'b0000010100100010;
            15'd19693: log10_cal = 16'b0000010100100010;
            15'd19694: log10_cal = 16'b0000010100100010;
            15'd19695: log10_cal = 16'b0000010100100010;
            15'd19696: log10_cal = 16'b0000010100100010;
            15'd19697: log10_cal = 16'b0000010100100010;
            15'd19698: log10_cal = 16'b0000010100100010;
            15'd19699: log10_cal = 16'b0000010100100010;
            15'd19700: log10_cal = 16'b0000010100100010;
            15'd19701: log10_cal = 16'b0000010100100011;
            15'd19702: log10_cal = 16'b0000010100100011;
            15'd19703: log10_cal = 16'b0000010100100011;
            15'd19704: log10_cal = 16'b0000010100100011;
            15'd19705: log10_cal = 16'b0000010100100011;
            15'd19706: log10_cal = 16'b0000010100100011;
            15'd19707: log10_cal = 16'b0000010100100011;
            15'd19708: log10_cal = 16'b0000010100100011;
            15'd19709: log10_cal = 16'b0000010100100011;
            15'd19710: log10_cal = 16'b0000010100100011;
            15'd19711: log10_cal = 16'b0000010100100011;
            15'd19712: log10_cal = 16'b0000010100100011;
            15'd19713: log10_cal = 16'b0000010100100011;
            15'd19714: log10_cal = 16'b0000010100100011;
            15'd19715: log10_cal = 16'b0000010100100011;
            15'd19716: log10_cal = 16'b0000010100100011;
            15'd19717: log10_cal = 16'b0000010100100011;
            15'd19718: log10_cal = 16'b0000010100100011;
            15'd19719: log10_cal = 16'b0000010100100011;
            15'd19720: log10_cal = 16'b0000010100100011;
            15'd19721: log10_cal = 16'b0000010100100011;
            15'd19722: log10_cal = 16'b0000010100100011;
            15'd19723: log10_cal = 16'b0000010100100011;
            15'd19724: log10_cal = 16'b0000010100100011;
            15'd19725: log10_cal = 16'b0000010100100011;
            15'd19726: log10_cal = 16'b0000010100100011;
            15'd19727: log10_cal = 16'b0000010100100011;
            15'd19728: log10_cal = 16'b0000010100100011;
            15'd19729: log10_cal = 16'b0000010100100011;
            15'd19730: log10_cal = 16'b0000010100100011;
            15'd19731: log10_cal = 16'b0000010100100011;
            15'd19732: log10_cal = 16'b0000010100100011;
            15'd19733: log10_cal = 16'b0000010100100011;
            15'd19734: log10_cal = 16'b0000010100100011;
            15'd19735: log10_cal = 16'b0000010100100011;
            15'd19736: log10_cal = 16'b0000010100100011;
            15'd19737: log10_cal = 16'b0000010100100011;
            15'd19738: log10_cal = 16'b0000010100100011;
            15'd19739: log10_cal = 16'b0000010100100011;
            15'd19740: log10_cal = 16'b0000010100100011;
            15'd19741: log10_cal = 16'b0000010100100011;
            15'd19742: log10_cal = 16'b0000010100100011;
            15'd19743: log10_cal = 16'b0000010100100011;
            15'd19744: log10_cal = 16'b0000010100100011;
            15'd19745: log10_cal = 16'b0000010100100100;
            15'd19746: log10_cal = 16'b0000010100100100;
            15'd19747: log10_cal = 16'b0000010100100100;
            15'd19748: log10_cal = 16'b0000010100100100;
            15'd19749: log10_cal = 16'b0000010100100100;
            15'd19750: log10_cal = 16'b0000010100100100;
            15'd19751: log10_cal = 16'b0000010100100100;
            15'd19752: log10_cal = 16'b0000010100100100;
            15'd19753: log10_cal = 16'b0000010100100100;
            15'd19754: log10_cal = 16'b0000010100100100;
            15'd19755: log10_cal = 16'b0000010100100100;
            15'd19756: log10_cal = 16'b0000010100100100;
            15'd19757: log10_cal = 16'b0000010100100100;
            15'd19758: log10_cal = 16'b0000010100100100;
            15'd19759: log10_cal = 16'b0000010100100100;
            15'd19760: log10_cal = 16'b0000010100100100;
            15'd19761: log10_cal = 16'b0000010100100100;
            15'd19762: log10_cal = 16'b0000010100100100;
            15'd19763: log10_cal = 16'b0000010100100100;
            15'd19764: log10_cal = 16'b0000010100100100;
            15'd19765: log10_cal = 16'b0000010100100100;
            15'd19766: log10_cal = 16'b0000010100100100;
            15'd19767: log10_cal = 16'b0000010100100100;
            15'd19768: log10_cal = 16'b0000010100100100;
            15'd19769: log10_cal = 16'b0000010100100100;
            15'd19770: log10_cal = 16'b0000010100100100;
            15'd19771: log10_cal = 16'b0000010100100100;
            15'd19772: log10_cal = 16'b0000010100100100;
            15'd19773: log10_cal = 16'b0000010100100100;
            15'd19774: log10_cal = 16'b0000010100100100;
            15'd19775: log10_cal = 16'b0000010100100100;
            15'd19776: log10_cal = 16'b0000010100100100;
            15'd19777: log10_cal = 16'b0000010100100100;
            15'd19778: log10_cal = 16'b0000010100100100;
            15'd19779: log10_cal = 16'b0000010100100100;
            15'd19780: log10_cal = 16'b0000010100100100;
            15'd19781: log10_cal = 16'b0000010100100100;
            15'd19782: log10_cal = 16'b0000010100100100;
            15'd19783: log10_cal = 16'b0000010100100100;
            15'd19784: log10_cal = 16'b0000010100100100;
            15'd19785: log10_cal = 16'b0000010100100100;
            15'd19786: log10_cal = 16'b0000010100100100;
            15'd19787: log10_cal = 16'b0000010100100100;
            15'd19788: log10_cal = 16'b0000010100100100;
            15'd19789: log10_cal = 16'b0000010100100100;
            15'd19790: log10_cal = 16'b0000010100100101;
            15'd19791: log10_cal = 16'b0000010100100101;
            15'd19792: log10_cal = 16'b0000010100100101;
            15'd19793: log10_cal = 16'b0000010100100101;
            15'd19794: log10_cal = 16'b0000010100100101;
            15'd19795: log10_cal = 16'b0000010100100101;
            15'd19796: log10_cal = 16'b0000010100100101;
            15'd19797: log10_cal = 16'b0000010100100101;
            15'd19798: log10_cal = 16'b0000010100100101;
            15'd19799: log10_cal = 16'b0000010100100101;
            15'd19800: log10_cal = 16'b0000010100100101;
            15'd19801: log10_cal = 16'b0000010100100101;
            15'd19802: log10_cal = 16'b0000010100100101;
            15'd19803: log10_cal = 16'b0000010100100101;
            15'd19804: log10_cal = 16'b0000010100100101;
            15'd19805: log10_cal = 16'b0000010100100101;
            15'd19806: log10_cal = 16'b0000010100100101;
            15'd19807: log10_cal = 16'b0000010100100101;
            15'd19808: log10_cal = 16'b0000010100100101;
            15'd19809: log10_cal = 16'b0000010100100101;
            15'd19810: log10_cal = 16'b0000010100100101;
            15'd19811: log10_cal = 16'b0000010100100101;
            15'd19812: log10_cal = 16'b0000010100100101;
            15'd19813: log10_cal = 16'b0000010100100101;
            15'd19814: log10_cal = 16'b0000010100100101;
            15'd19815: log10_cal = 16'b0000010100100101;
            15'd19816: log10_cal = 16'b0000010100100101;
            15'd19817: log10_cal = 16'b0000010100100101;
            15'd19818: log10_cal = 16'b0000010100100101;
            15'd19819: log10_cal = 16'b0000010100100101;
            15'd19820: log10_cal = 16'b0000010100100101;
            15'd19821: log10_cal = 16'b0000010100100101;
            15'd19822: log10_cal = 16'b0000010100100101;
            15'd19823: log10_cal = 16'b0000010100100101;
            15'd19824: log10_cal = 16'b0000010100100101;
            15'd19825: log10_cal = 16'b0000010100100101;
            15'd19826: log10_cal = 16'b0000010100100101;
            15'd19827: log10_cal = 16'b0000010100100101;
            15'd19828: log10_cal = 16'b0000010100100101;
            15'd19829: log10_cal = 16'b0000010100100101;
            15'd19830: log10_cal = 16'b0000010100100101;
            15'd19831: log10_cal = 16'b0000010100100101;
            15'd19832: log10_cal = 16'b0000010100100101;
            15'd19833: log10_cal = 16'b0000010100100101;
            15'd19834: log10_cal = 16'b0000010100100110;
            15'd19835: log10_cal = 16'b0000010100100110;
            15'd19836: log10_cal = 16'b0000010100100110;
            15'd19837: log10_cal = 16'b0000010100100110;
            15'd19838: log10_cal = 16'b0000010100100110;
            15'd19839: log10_cal = 16'b0000010100100110;
            15'd19840: log10_cal = 16'b0000010100100110;
            15'd19841: log10_cal = 16'b0000010100100110;
            15'd19842: log10_cal = 16'b0000010100100110;
            15'd19843: log10_cal = 16'b0000010100100110;
            15'd19844: log10_cal = 16'b0000010100100110;
            15'd19845: log10_cal = 16'b0000010100100110;
            15'd19846: log10_cal = 16'b0000010100100110;
            15'd19847: log10_cal = 16'b0000010100100110;
            15'd19848: log10_cal = 16'b0000010100100110;
            15'd19849: log10_cal = 16'b0000010100100110;
            15'd19850: log10_cal = 16'b0000010100100110;
            15'd19851: log10_cal = 16'b0000010100100110;
            15'd19852: log10_cal = 16'b0000010100100110;
            15'd19853: log10_cal = 16'b0000010100100110;
            15'd19854: log10_cal = 16'b0000010100100110;
            15'd19855: log10_cal = 16'b0000010100100110;
            15'd19856: log10_cal = 16'b0000010100100110;
            15'd19857: log10_cal = 16'b0000010100100110;
            15'd19858: log10_cal = 16'b0000010100100110;
            15'd19859: log10_cal = 16'b0000010100100110;
            15'd19860: log10_cal = 16'b0000010100100110;
            15'd19861: log10_cal = 16'b0000010100100110;
            15'd19862: log10_cal = 16'b0000010100100110;
            15'd19863: log10_cal = 16'b0000010100100110;
            15'd19864: log10_cal = 16'b0000010100100110;
            15'd19865: log10_cal = 16'b0000010100100110;
            15'd19866: log10_cal = 16'b0000010100100110;
            15'd19867: log10_cal = 16'b0000010100100110;
            15'd19868: log10_cal = 16'b0000010100100110;
            15'd19869: log10_cal = 16'b0000010100100110;
            15'd19870: log10_cal = 16'b0000010100100110;
            15'd19871: log10_cal = 16'b0000010100100110;
            15'd19872: log10_cal = 16'b0000010100100110;
            15'd19873: log10_cal = 16'b0000010100100110;
            15'd19874: log10_cal = 16'b0000010100100110;
            15'd19875: log10_cal = 16'b0000010100100110;
            15'd19876: log10_cal = 16'b0000010100100110;
            15'd19877: log10_cal = 16'b0000010100100110;
            15'd19878: log10_cal = 16'b0000010100100110;
            15'd19879: log10_cal = 16'b0000010100100111;
            15'd19880: log10_cal = 16'b0000010100100111;
            15'd19881: log10_cal = 16'b0000010100100111;
            15'd19882: log10_cal = 16'b0000010100100111;
            15'd19883: log10_cal = 16'b0000010100100111;
            15'd19884: log10_cal = 16'b0000010100100111;
            15'd19885: log10_cal = 16'b0000010100100111;
            15'd19886: log10_cal = 16'b0000010100100111;
            15'd19887: log10_cal = 16'b0000010100100111;
            15'd19888: log10_cal = 16'b0000010100100111;
            15'd19889: log10_cal = 16'b0000010100100111;
            15'd19890: log10_cal = 16'b0000010100100111;
            15'd19891: log10_cal = 16'b0000010100100111;
            15'd19892: log10_cal = 16'b0000010100100111;
            15'd19893: log10_cal = 16'b0000010100100111;
            15'd19894: log10_cal = 16'b0000010100100111;
            15'd19895: log10_cal = 16'b0000010100100111;
            15'd19896: log10_cal = 16'b0000010100100111;
            15'd19897: log10_cal = 16'b0000010100100111;
            15'd19898: log10_cal = 16'b0000010100100111;
            15'd19899: log10_cal = 16'b0000010100100111;
            15'd19900: log10_cal = 16'b0000010100100111;
            15'd19901: log10_cal = 16'b0000010100100111;
            15'd19902: log10_cal = 16'b0000010100100111;
            15'd19903: log10_cal = 16'b0000010100100111;
            15'd19904: log10_cal = 16'b0000010100100111;
            15'd19905: log10_cal = 16'b0000010100100111;
            15'd19906: log10_cal = 16'b0000010100100111;
            15'd19907: log10_cal = 16'b0000010100100111;
            15'd19908: log10_cal = 16'b0000010100100111;
            15'd19909: log10_cal = 16'b0000010100100111;
            15'd19910: log10_cal = 16'b0000010100100111;
            15'd19911: log10_cal = 16'b0000010100100111;
            15'd19912: log10_cal = 16'b0000010100100111;
            15'd19913: log10_cal = 16'b0000010100100111;
            15'd19914: log10_cal = 16'b0000010100100111;
            15'd19915: log10_cal = 16'b0000010100100111;
            15'd19916: log10_cal = 16'b0000010100100111;
            15'd19917: log10_cal = 16'b0000010100100111;
            15'd19918: log10_cal = 16'b0000010100100111;
            15'd19919: log10_cal = 16'b0000010100100111;
            15'd19920: log10_cal = 16'b0000010100100111;
            15'd19921: log10_cal = 16'b0000010100100111;
            15'd19922: log10_cal = 16'b0000010100100111;
            15'd19923: log10_cal = 16'b0000010100100111;
            15'd19924: log10_cal = 16'b0000010100101000;
            15'd19925: log10_cal = 16'b0000010100101000;
            15'd19926: log10_cal = 16'b0000010100101000;
            15'd19927: log10_cal = 16'b0000010100101000;
            15'd19928: log10_cal = 16'b0000010100101000;
            15'd19929: log10_cal = 16'b0000010100101000;
            15'd19930: log10_cal = 16'b0000010100101000;
            15'd19931: log10_cal = 16'b0000010100101000;
            15'd19932: log10_cal = 16'b0000010100101000;
            15'd19933: log10_cal = 16'b0000010100101000;
            15'd19934: log10_cal = 16'b0000010100101000;
            15'd19935: log10_cal = 16'b0000010100101000;
            15'd19936: log10_cal = 16'b0000010100101000;
            15'd19937: log10_cal = 16'b0000010100101000;
            15'd19938: log10_cal = 16'b0000010100101000;
            15'd19939: log10_cal = 16'b0000010100101000;
            15'd19940: log10_cal = 16'b0000010100101000;
            15'd19941: log10_cal = 16'b0000010100101000;
            15'd19942: log10_cal = 16'b0000010100101000;
            15'd19943: log10_cal = 16'b0000010100101000;
            15'd19944: log10_cal = 16'b0000010100101000;
            15'd19945: log10_cal = 16'b0000010100101000;
            15'd19946: log10_cal = 16'b0000010100101000;
            15'd19947: log10_cal = 16'b0000010100101000;
            15'd19948: log10_cal = 16'b0000010100101000;
            15'd19949: log10_cal = 16'b0000010100101000;
            15'd19950: log10_cal = 16'b0000010100101000;
            15'd19951: log10_cal = 16'b0000010100101000;
            15'd19952: log10_cal = 16'b0000010100101000;
            15'd19953: log10_cal = 16'b0000010100101000;
            15'd19954: log10_cal = 16'b0000010100101000;
            15'd19955: log10_cal = 16'b0000010100101000;
            15'd19956: log10_cal = 16'b0000010100101000;
            15'd19957: log10_cal = 16'b0000010100101000;
            15'd19958: log10_cal = 16'b0000010100101000;
            15'd19959: log10_cal = 16'b0000010100101000;
            15'd19960: log10_cal = 16'b0000010100101000;
            15'd19961: log10_cal = 16'b0000010100101000;
            15'd19962: log10_cal = 16'b0000010100101000;
            15'd19963: log10_cal = 16'b0000010100101000;
            15'd19964: log10_cal = 16'b0000010100101000;
            15'd19965: log10_cal = 16'b0000010100101000;
            15'd19966: log10_cal = 16'b0000010100101000;
            15'd19967: log10_cal = 16'b0000010100101000;
            15'd19968: log10_cal = 16'b0000010100101000;
            15'd19969: log10_cal = 16'b0000010100101001;
            15'd19970: log10_cal = 16'b0000010100101001;
            15'd19971: log10_cal = 16'b0000010100101001;
            15'd19972: log10_cal = 16'b0000010100101001;
            15'd19973: log10_cal = 16'b0000010100101001;
            15'd19974: log10_cal = 16'b0000010100101001;
            15'd19975: log10_cal = 16'b0000010100101001;
            15'd19976: log10_cal = 16'b0000010100101001;
            15'd19977: log10_cal = 16'b0000010100101001;
            15'd19978: log10_cal = 16'b0000010100101001;
            15'd19979: log10_cal = 16'b0000010100101001;
            15'd19980: log10_cal = 16'b0000010100101001;
            15'd19981: log10_cal = 16'b0000010100101001;
            15'd19982: log10_cal = 16'b0000010100101001;
            15'd19983: log10_cal = 16'b0000010100101001;
            15'd19984: log10_cal = 16'b0000010100101001;
            15'd19985: log10_cal = 16'b0000010100101001;
            15'd19986: log10_cal = 16'b0000010100101001;
            15'd19987: log10_cal = 16'b0000010100101001;
            15'd19988: log10_cal = 16'b0000010100101001;
            15'd19989: log10_cal = 16'b0000010100101001;
            15'd19990: log10_cal = 16'b0000010100101001;
            15'd19991: log10_cal = 16'b0000010100101001;
            15'd19992: log10_cal = 16'b0000010100101001;
            15'd19993: log10_cal = 16'b0000010100101001;
            15'd19994: log10_cal = 16'b0000010100101001;
            15'd19995: log10_cal = 16'b0000010100101001;
            15'd19996: log10_cal = 16'b0000010100101001;
            15'd19997: log10_cal = 16'b0000010100101001;
            15'd19998: log10_cal = 16'b0000010100101001;
            15'd19999: log10_cal = 16'b0000010100101001;
            15'd20000: log10_cal = 16'b0000010100101001;
            15'd20001: log10_cal = 16'b0000010100101001;
            15'd20002: log10_cal = 16'b0000010100101001;
            15'd20003: log10_cal = 16'b0000010100101001;
            15'd20004: log10_cal = 16'b0000010100101001;
            15'd20005: log10_cal = 16'b0000010100101001;
            15'd20006: log10_cal = 16'b0000010100101001;
            15'd20007: log10_cal = 16'b0000010100101001;
            15'd20008: log10_cal = 16'b0000010100101001;
            15'd20009: log10_cal = 16'b0000010100101001;
            15'd20010: log10_cal = 16'b0000010100101001;
            15'd20011: log10_cal = 16'b0000010100101001;
            15'd20012: log10_cal = 16'b0000010100101001;
            15'd20013: log10_cal = 16'b0000010100101001;
            15'd20014: log10_cal = 16'b0000010100101010;
            15'd20015: log10_cal = 16'b0000010100101010;
            15'd20016: log10_cal = 16'b0000010100101010;
            15'd20017: log10_cal = 16'b0000010100101010;
            15'd20018: log10_cal = 16'b0000010100101010;
            15'd20019: log10_cal = 16'b0000010100101010;
            15'd20020: log10_cal = 16'b0000010100101010;
            15'd20021: log10_cal = 16'b0000010100101010;
            15'd20022: log10_cal = 16'b0000010100101010;
            15'd20023: log10_cal = 16'b0000010100101010;
            15'd20024: log10_cal = 16'b0000010100101010;
            15'd20025: log10_cal = 16'b0000010100101010;
            15'd20026: log10_cal = 16'b0000010100101010;
            15'd20027: log10_cal = 16'b0000010100101010;
            15'd20028: log10_cal = 16'b0000010100101010;
            15'd20029: log10_cal = 16'b0000010100101010;
            15'd20030: log10_cal = 16'b0000010100101010;
            15'd20031: log10_cal = 16'b0000010100101010;
            15'd20032: log10_cal = 16'b0000010100101010;
            15'd20033: log10_cal = 16'b0000010100101010;
            15'd20034: log10_cal = 16'b0000010100101010;
            15'd20035: log10_cal = 16'b0000010100101010;
            15'd20036: log10_cal = 16'b0000010100101010;
            15'd20037: log10_cal = 16'b0000010100101010;
            15'd20038: log10_cal = 16'b0000010100101010;
            15'd20039: log10_cal = 16'b0000010100101010;
            15'd20040: log10_cal = 16'b0000010100101010;
            15'd20041: log10_cal = 16'b0000010100101010;
            15'd20042: log10_cal = 16'b0000010100101010;
            15'd20043: log10_cal = 16'b0000010100101010;
            15'd20044: log10_cal = 16'b0000010100101010;
            15'd20045: log10_cal = 16'b0000010100101010;
            15'd20046: log10_cal = 16'b0000010100101010;
            15'd20047: log10_cal = 16'b0000010100101010;
            15'd20048: log10_cal = 16'b0000010100101010;
            15'd20049: log10_cal = 16'b0000010100101010;
            15'd20050: log10_cal = 16'b0000010100101010;
            15'd20051: log10_cal = 16'b0000010100101010;
            15'd20052: log10_cal = 16'b0000010100101010;
            15'd20053: log10_cal = 16'b0000010100101010;
            15'd20054: log10_cal = 16'b0000010100101010;
            15'd20055: log10_cal = 16'b0000010100101010;
            15'd20056: log10_cal = 16'b0000010100101010;
            15'd20057: log10_cal = 16'b0000010100101010;
            15'd20058: log10_cal = 16'b0000010100101010;
            15'd20059: log10_cal = 16'b0000010100101011;
            15'd20060: log10_cal = 16'b0000010100101011;
            15'd20061: log10_cal = 16'b0000010100101011;
            15'd20062: log10_cal = 16'b0000010100101011;
            15'd20063: log10_cal = 16'b0000010100101011;
            15'd20064: log10_cal = 16'b0000010100101011;
            15'd20065: log10_cal = 16'b0000010100101011;
            15'd20066: log10_cal = 16'b0000010100101011;
            15'd20067: log10_cal = 16'b0000010100101011;
            15'd20068: log10_cal = 16'b0000010100101011;
            15'd20069: log10_cal = 16'b0000010100101011;
            15'd20070: log10_cal = 16'b0000010100101011;
            15'd20071: log10_cal = 16'b0000010100101011;
            15'd20072: log10_cal = 16'b0000010100101011;
            15'd20073: log10_cal = 16'b0000010100101011;
            15'd20074: log10_cal = 16'b0000010100101011;
            15'd20075: log10_cal = 16'b0000010100101011;
            15'd20076: log10_cal = 16'b0000010100101011;
            15'd20077: log10_cal = 16'b0000010100101011;
            15'd20078: log10_cal = 16'b0000010100101011;
            15'd20079: log10_cal = 16'b0000010100101011;
            15'd20080: log10_cal = 16'b0000010100101011;
            15'd20081: log10_cal = 16'b0000010100101011;
            15'd20082: log10_cal = 16'b0000010100101011;
            15'd20083: log10_cal = 16'b0000010100101011;
            15'd20084: log10_cal = 16'b0000010100101011;
            15'd20085: log10_cal = 16'b0000010100101011;
            15'd20086: log10_cal = 16'b0000010100101011;
            15'd20087: log10_cal = 16'b0000010100101011;
            15'd20088: log10_cal = 16'b0000010100101011;
            15'd20089: log10_cal = 16'b0000010100101011;
            15'd20090: log10_cal = 16'b0000010100101011;
            15'd20091: log10_cal = 16'b0000010100101011;
            15'd20092: log10_cal = 16'b0000010100101011;
            15'd20093: log10_cal = 16'b0000010100101011;
            15'd20094: log10_cal = 16'b0000010100101011;
            15'd20095: log10_cal = 16'b0000010100101011;
            15'd20096: log10_cal = 16'b0000010100101011;
            15'd20097: log10_cal = 16'b0000010100101011;
            15'd20098: log10_cal = 16'b0000010100101011;
            15'd20099: log10_cal = 16'b0000010100101011;
            15'd20100: log10_cal = 16'b0000010100101011;
            15'd20101: log10_cal = 16'b0000010100101011;
            15'd20102: log10_cal = 16'b0000010100101011;
            15'd20103: log10_cal = 16'b0000010100101011;
            15'd20104: log10_cal = 16'b0000010100101100;
            15'd20105: log10_cal = 16'b0000010100101100;
            15'd20106: log10_cal = 16'b0000010100101100;
            15'd20107: log10_cal = 16'b0000010100101100;
            15'd20108: log10_cal = 16'b0000010100101100;
            15'd20109: log10_cal = 16'b0000010100101100;
            15'd20110: log10_cal = 16'b0000010100101100;
            15'd20111: log10_cal = 16'b0000010100101100;
            15'd20112: log10_cal = 16'b0000010100101100;
            15'd20113: log10_cal = 16'b0000010100101100;
            15'd20114: log10_cal = 16'b0000010100101100;
            15'd20115: log10_cal = 16'b0000010100101100;
            15'd20116: log10_cal = 16'b0000010100101100;
            15'd20117: log10_cal = 16'b0000010100101100;
            15'd20118: log10_cal = 16'b0000010100101100;
            15'd20119: log10_cal = 16'b0000010100101100;
            15'd20120: log10_cal = 16'b0000010100101100;
            15'd20121: log10_cal = 16'b0000010100101100;
            15'd20122: log10_cal = 16'b0000010100101100;
            15'd20123: log10_cal = 16'b0000010100101100;
            15'd20124: log10_cal = 16'b0000010100101100;
            15'd20125: log10_cal = 16'b0000010100101100;
            15'd20126: log10_cal = 16'b0000010100101100;
            15'd20127: log10_cal = 16'b0000010100101100;
            15'd20128: log10_cal = 16'b0000010100101100;
            15'd20129: log10_cal = 16'b0000010100101100;
            15'd20130: log10_cal = 16'b0000010100101100;
            15'd20131: log10_cal = 16'b0000010100101100;
            15'd20132: log10_cal = 16'b0000010100101100;
            15'd20133: log10_cal = 16'b0000010100101100;
            15'd20134: log10_cal = 16'b0000010100101100;
            15'd20135: log10_cal = 16'b0000010100101100;
            15'd20136: log10_cal = 16'b0000010100101100;
            15'd20137: log10_cal = 16'b0000010100101100;
            15'd20138: log10_cal = 16'b0000010100101100;
            15'd20139: log10_cal = 16'b0000010100101100;
            15'd20140: log10_cal = 16'b0000010100101100;
            15'd20141: log10_cal = 16'b0000010100101100;
            15'd20142: log10_cal = 16'b0000010100101100;
            15'd20143: log10_cal = 16'b0000010100101100;
            15'd20144: log10_cal = 16'b0000010100101100;
            15'd20145: log10_cal = 16'b0000010100101100;
            15'd20146: log10_cal = 16'b0000010100101100;
            15'd20147: log10_cal = 16'b0000010100101100;
            15'd20148: log10_cal = 16'b0000010100101100;
            15'd20149: log10_cal = 16'b0000010100101101;
            15'd20150: log10_cal = 16'b0000010100101101;
            15'd20151: log10_cal = 16'b0000010100101101;
            15'd20152: log10_cal = 16'b0000010100101101;
            15'd20153: log10_cal = 16'b0000010100101101;
            15'd20154: log10_cal = 16'b0000010100101101;
            15'd20155: log10_cal = 16'b0000010100101101;
            15'd20156: log10_cal = 16'b0000010100101101;
            15'd20157: log10_cal = 16'b0000010100101101;
            15'd20158: log10_cal = 16'b0000010100101101;
            15'd20159: log10_cal = 16'b0000010100101101;
            15'd20160: log10_cal = 16'b0000010100101101;
            15'd20161: log10_cal = 16'b0000010100101101;
            15'd20162: log10_cal = 16'b0000010100101101;
            15'd20163: log10_cal = 16'b0000010100101101;
            15'd20164: log10_cal = 16'b0000010100101101;
            15'd20165: log10_cal = 16'b0000010100101101;
            15'd20166: log10_cal = 16'b0000010100101101;
            15'd20167: log10_cal = 16'b0000010100101101;
            15'd20168: log10_cal = 16'b0000010100101101;
            15'd20169: log10_cal = 16'b0000010100101101;
            15'd20170: log10_cal = 16'b0000010100101101;
            15'd20171: log10_cal = 16'b0000010100101101;
            15'd20172: log10_cal = 16'b0000010100101101;
            15'd20173: log10_cal = 16'b0000010100101101;
            15'd20174: log10_cal = 16'b0000010100101101;
            15'd20175: log10_cal = 16'b0000010100101101;
            15'd20176: log10_cal = 16'b0000010100101101;
            15'd20177: log10_cal = 16'b0000010100101101;
            15'd20178: log10_cal = 16'b0000010100101101;
            15'd20179: log10_cal = 16'b0000010100101101;
            15'd20180: log10_cal = 16'b0000010100101101;
            15'd20181: log10_cal = 16'b0000010100101101;
            15'd20182: log10_cal = 16'b0000010100101101;
            15'd20183: log10_cal = 16'b0000010100101101;
            15'd20184: log10_cal = 16'b0000010100101101;
            15'd20185: log10_cal = 16'b0000010100101101;
            15'd20186: log10_cal = 16'b0000010100101101;
            15'd20187: log10_cal = 16'b0000010100101101;
            15'd20188: log10_cal = 16'b0000010100101101;
            15'd20189: log10_cal = 16'b0000010100101101;
            15'd20190: log10_cal = 16'b0000010100101101;
            15'd20191: log10_cal = 16'b0000010100101101;
            15'd20192: log10_cal = 16'b0000010100101101;
            15'd20193: log10_cal = 16'b0000010100101101;
            15'd20194: log10_cal = 16'b0000010100101110;
            15'd20195: log10_cal = 16'b0000010100101110;
            15'd20196: log10_cal = 16'b0000010100101110;
            15'd20197: log10_cal = 16'b0000010100101110;
            15'd20198: log10_cal = 16'b0000010100101110;
            15'd20199: log10_cal = 16'b0000010100101110;
            15'd20200: log10_cal = 16'b0000010100101110;
            15'd20201: log10_cal = 16'b0000010100101110;
            15'd20202: log10_cal = 16'b0000010100101110;
            15'd20203: log10_cal = 16'b0000010100101110;
            15'd20204: log10_cal = 16'b0000010100101110;
            15'd20205: log10_cal = 16'b0000010100101110;
            15'd20206: log10_cal = 16'b0000010100101110;
            15'd20207: log10_cal = 16'b0000010100101110;
            15'd20208: log10_cal = 16'b0000010100101110;
            15'd20209: log10_cal = 16'b0000010100101110;
            15'd20210: log10_cal = 16'b0000010100101110;
            15'd20211: log10_cal = 16'b0000010100101110;
            15'd20212: log10_cal = 16'b0000010100101110;
            15'd20213: log10_cal = 16'b0000010100101110;
            15'd20214: log10_cal = 16'b0000010100101110;
            15'd20215: log10_cal = 16'b0000010100101110;
            15'd20216: log10_cal = 16'b0000010100101110;
            15'd20217: log10_cal = 16'b0000010100101110;
            15'd20218: log10_cal = 16'b0000010100101110;
            15'd20219: log10_cal = 16'b0000010100101110;
            15'd20220: log10_cal = 16'b0000010100101110;
            15'd20221: log10_cal = 16'b0000010100101110;
            15'd20222: log10_cal = 16'b0000010100101110;
            15'd20223: log10_cal = 16'b0000010100101110;
            15'd20224: log10_cal = 16'b0000010100101110;
            15'd20225: log10_cal = 16'b0000010100101110;
            15'd20226: log10_cal = 16'b0000010100101110;
            15'd20227: log10_cal = 16'b0000010100101110;
            15'd20228: log10_cal = 16'b0000010100101110;
            15'd20229: log10_cal = 16'b0000010100101110;
            15'd20230: log10_cal = 16'b0000010100101110;
            15'd20231: log10_cal = 16'b0000010100101110;
            15'd20232: log10_cal = 16'b0000010100101110;
            15'd20233: log10_cal = 16'b0000010100101110;
            15'd20234: log10_cal = 16'b0000010100101110;
            15'd20235: log10_cal = 16'b0000010100101110;
            15'd20236: log10_cal = 16'b0000010100101110;
            15'd20237: log10_cal = 16'b0000010100101110;
            15'd20238: log10_cal = 16'b0000010100101110;
            15'd20239: log10_cal = 16'b0000010100101110;
            15'd20240: log10_cal = 16'b0000010100101111;
            15'd20241: log10_cal = 16'b0000010100101111;
            15'd20242: log10_cal = 16'b0000010100101111;
            15'd20243: log10_cal = 16'b0000010100101111;
            15'd20244: log10_cal = 16'b0000010100101111;
            15'd20245: log10_cal = 16'b0000010100101111;
            15'd20246: log10_cal = 16'b0000010100101111;
            15'd20247: log10_cal = 16'b0000010100101111;
            15'd20248: log10_cal = 16'b0000010100101111;
            15'd20249: log10_cal = 16'b0000010100101111;
            15'd20250: log10_cal = 16'b0000010100101111;
            15'd20251: log10_cal = 16'b0000010100101111;
            15'd20252: log10_cal = 16'b0000010100101111;
            15'd20253: log10_cal = 16'b0000010100101111;
            15'd20254: log10_cal = 16'b0000010100101111;
            15'd20255: log10_cal = 16'b0000010100101111;
            15'd20256: log10_cal = 16'b0000010100101111;
            15'd20257: log10_cal = 16'b0000010100101111;
            15'd20258: log10_cal = 16'b0000010100101111;
            15'd20259: log10_cal = 16'b0000010100101111;
            15'd20260: log10_cal = 16'b0000010100101111;
            15'd20261: log10_cal = 16'b0000010100101111;
            15'd20262: log10_cal = 16'b0000010100101111;
            15'd20263: log10_cal = 16'b0000010100101111;
            15'd20264: log10_cal = 16'b0000010100101111;
            15'd20265: log10_cal = 16'b0000010100101111;
            15'd20266: log10_cal = 16'b0000010100101111;
            15'd20267: log10_cal = 16'b0000010100101111;
            15'd20268: log10_cal = 16'b0000010100101111;
            15'd20269: log10_cal = 16'b0000010100101111;
            15'd20270: log10_cal = 16'b0000010100101111;
            15'd20271: log10_cal = 16'b0000010100101111;
            15'd20272: log10_cal = 16'b0000010100101111;
            15'd20273: log10_cal = 16'b0000010100101111;
            15'd20274: log10_cal = 16'b0000010100101111;
            15'd20275: log10_cal = 16'b0000010100101111;
            15'd20276: log10_cal = 16'b0000010100101111;
            15'd20277: log10_cal = 16'b0000010100101111;
            15'd20278: log10_cal = 16'b0000010100101111;
            15'd20279: log10_cal = 16'b0000010100101111;
            15'd20280: log10_cal = 16'b0000010100101111;
            15'd20281: log10_cal = 16'b0000010100101111;
            15'd20282: log10_cal = 16'b0000010100101111;
            15'd20283: log10_cal = 16'b0000010100101111;
            15'd20284: log10_cal = 16'b0000010100101111;
            15'd20285: log10_cal = 16'b0000010100110000;
            15'd20286: log10_cal = 16'b0000010100110000;
            15'd20287: log10_cal = 16'b0000010100110000;
            15'd20288: log10_cal = 16'b0000010100110000;
            15'd20289: log10_cal = 16'b0000010100110000;
            15'd20290: log10_cal = 16'b0000010100110000;
            15'd20291: log10_cal = 16'b0000010100110000;
            15'd20292: log10_cal = 16'b0000010100110000;
            15'd20293: log10_cal = 16'b0000010100110000;
            15'd20294: log10_cal = 16'b0000010100110000;
            15'd20295: log10_cal = 16'b0000010100110000;
            15'd20296: log10_cal = 16'b0000010100110000;
            15'd20297: log10_cal = 16'b0000010100110000;
            15'd20298: log10_cal = 16'b0000010100110000;
            15'd20299: log10_cal = 16'b0000010100110000;
            15'd20300: log10_cal = 16'b0000010100110000;
            15'd20301: log10_cal = 16'b0000010100110000;
            15'd20302: log10_cal = 16'b0000010100110000;
            15'd20303: log10_cal = 16'b0000010100110000;
            15'd20304: log10_cal = 16'b0000010100110000;
            15'd20305: log10_cal = 16'b0000010100110000;
            15'd20306: log10_cal = 16'b0000010100110000;
            15'd20307: log10_cal = 16'b0000010100110000;
            15'd20308: log10_cal = 16'b0000010100110000;
            15'd20309: log10_cal = 16'b0000010100110000;
            15'd20310: log10_cal = 16'b0000010100110000;
            15'd20311: log10_cal = 16'b0000010100110000;
            15'd20312: log10_cal = 16'b0000010100110000;
            15'd20313: log10_cal = 16'b0000010100110000;
            15'd20314: log10_cal = 16'b0000010100110000;
            15'd20315: log10_cal = 16'b0000010100110000;
            15'd20316: log10_cal = 16'b0000010100110000;
            15'd20317: log10_cal = 16'b0000010100110000;
            15'd20318: log10_cal = 16'b0000010100110000;
            15'd20319: log10_cal = 16'b0000010100110000;
            15'd20320: log10_cal = 16'b0000010100110000;
            15'd20321: log10_cal = 16'b0000010100110000;
            15'd20322: log10_cal = 16'b0000010100110000;
            15'd20323: log10_cal = 16'b0000010100110000;
            15'd20324: log10_cal = 16'b0000010100110000;
            15'd20325: log10_cal = 16'b0000010100110000;
            15'd20326: log10_cal = 16'b0000010100110000;
            15'd20327: log10_cal = 16'b0000010100110000;
            15'd20328: log10_cal = 16'b0000010100110000;
            15'd20329: log10_cal = 16'b0000010100110000;
            15'd20330: log10_cal = 16'b0000010100110000;
            15'd20331: log10_cal = 16'b0000010100110001;
            15'd20332: log10_cal = 16'b0000010100110001;
            15'd20333: log10_cal = 16'b0000010100110001;
            15'd20334: log10_cal = 16'b0000010100110001;
            15'd20335: log10_cal = 16'b0000010100110001;
            15'd20336: log10_cal = 16'b0000010100110001;
            15'd20337: log10_cal = 16'b0000010100110001;
            15'd20338: log10_cal = 16'b0000010100110001;
            15'd20339: log10_cal = 16'b0000010100110001;
            15'd20340: log10_cal = 16'b0000010100110001;
            15'd20341: log10_cal = 16'b0000010100110001;
            15'd20342: log10_cal = 16'b0000010100110001;
            15'd20343: log10_cal = 16'b0000010100110001;
            15'd20344: log10_cal = 16'b0000010100110001;
            15'd20345: log10_cal = 16'b0000010100110001;
            15'd20346: log10_cal = 16'b0000010100110001;
            15'd20347: log10_cal = 16'b0000010100110001;
            15'd20348: log10_cal = 16'b0000010100110001;
            15'd20349: log10_cal = 16'b0000010100110001;
            15'd20350: log10_cal = 16'b0000010100110001;
            15'd20351: log10_cal = 16'b0000010100110001;
            15'd20352: log10_cal = 16'b0000010100110001;
            15'd20353: log10_cal = 16'b0000010100110001;
            15'd20354: log10_cal = 16'b0000010100110001;
            15'd20355: log10_cal = 16'b0000010100110001;
            15'd20356: log10_cal = 16'b0000010100110001;
            15'd20357: log10_cal = 16'b0000010100110001;
            15'd20358: log10_cal = 16'b0000010100110001;
            15'd20359: log10_cal = 16'b0000010100110001;
            15'd20360: log10_cal = 16'b0000010100110001;
            15'd20361: log10_cal = 16'b0000010100110001;
            15'd20362: log10_cal = 16'b0000010100110001;
            15'd20363: log10_cal = 16'b0000010100110001;
            15'd20364: log10_cal = 16'b0000010100110001;
            15'd20365: log10_cal = 16'b0000010100110001;
            15'd20366: log10_cal = 16'b0000010100110001;
            15'd20367: log10_cal = 16'b0000010100110001;
            15'd20368: log10_cal = 16'b0000010100110001;
            15'd20369: log10_cal = 16'b0000010100110001;
            15'd20370: log10_cal = 16'b0000010100110001;
            15'd20371: log10_cal = 16'b0000010100110001;
            15'd20372: log10_cal = 16'b0000010100110001;
            15'd20373: log10_cal = 16'b0000010100110001;
            15'd20374: log10_cal = 16'b0000010100110001;
            15'd20375: log10_cal = 16'b0000010100110001;
            15'd20376: log10_cal = 16'b0000010100110001;
            15'd20377: log10_cal = 16'b0000010100110010;
            15'd20378: log10_cal = 16'b0000010100110010;
            15'd20379: log10_cal = 16'b0000010100110010;
            15'd20380: log10_cal = 16'b0000010100110010;
            15'd20381: log10_cal = 16'b0000010100110010;
            15'd20382: log10_cal = 16'b0000010100110010;
            15'd20383: log10_cal = 16'b0000010100110010;
            15'd20384: log10_cal = 16'b0000010100110010;
            15'd20385: log10_cal = 16'b0000010100110010;
            15'd20386: log10_cal = 16'b0000010100110010;
            15'd20387: log10_cal = 16'b0000010100110010;
            15'd20388: log10_cal = 16'b0000010100110010;
            15'd20389: log10_cal = 16'b0000010100110010;
            15'd20390: log10_cal = 16'b0000010100110010;
            15'd20391: log10_cal = 16'b0000010100110010;
            15'd20392: log10_cal = 16'b0000010100110010;
            15'd20393: log10_cal = 16'b0000010100110010;
            15'd20394: log10_cal = 16'b0000010100110010;
            15'd20395: log10_cal = 16'b0000010100110010;
            15'd20396: log10_cal = 16'b0000010100110010;
            15'd20397: log10_cal = 16'b0000010100110010;
            15'd20398: log10_cal = 16'b0000010100110010;
            15'd20399: log10_cal = 16'b0000010100110010;
            15'd20400: log10_cal = 16'b0000010100110010;
            15'd20401: log10_cal = 16'b0000010100110010;
            15'd20402: log10_cal = 16'b0000010100110010;
            15'd20403: log10_cal = 16'b0000010100110010;
            15'd20404: log10_cal = 16'b0000010100110010;
            15'd20405: log10_cal = 16'b0000010100110010;
            15'd20406: log10_cal = 16'b0000010100110010;
            15'd20407: log10_cal = 16'b0000010100110010;
            15'd20408: log10_cal = 16'b0000010100110010;
            15'd20409: log10_cal = 16'b0000010100110010;
            15'd20410: log10_cal = 16'b0000010100110010;
            15'd20411: log10_cal = 16'b0000010100110010;
            15'd20412: log10_cal = 16'b0000010100110010;
            15'd20413: log10_cal = 16'b0000010100110010;
            15'd20414: log10_cal = 16'b0000010100110010;
            15'd20415: log10_cal = 16'b0000010100110010;
            15'd20416: log10_cal = 16'b0000010100110010;
            15'd20417: log10_cal = 16'b0000010100110010;
            15'd20418: log10_cal = 16'b0000010100110010;
            15'd20419: log10_cal = 16'b0000010100110010;
            15'd20420: log10_cal = 16'b0000010100110010;
            15'd20421: log10_cal = 16'b0000010100110010;
            15'd20422: log10_cal = 16'b0000010100110010;
            15'd20423: log10_cal = 16'b0000010100110011;
            15'd20424: log10_cal = 16'b0000010100110011;
            15'd20425: log10_cal = 16'b0000010100110011;
            15'd20426: log10_cal = 16'b0000010100110011;
            15'd20427: log10_cal = 16'b0000010100110011;
            15'd20428: log10_cal = 16'b0000010100110011;
            15'd20429: log10_cal = 16'b0000010100110011;
            15'd20430: log10_cal = 16'b0000010100110011;
            15'd20431: log10_cal = 16'b0000010100110011;
            15'd20432: log10_cal = 16'b0000010100110011;
            15'd20433: log10_cal = 16'b0000010100110011;
            15'd20434: log10_cal = 16'b0000010100110011;
            15'd20435: log10_cal = 16'b0000010100110011;
            15'd20436: log10_cal = 16'b0000010100110011;
            15'd20437: log10_cal = 16'b0000010100110011;
            15'd20438: log10_cal = 16'b0000010100110011;
            15'd20439: log10_cal = 16'b0000010100110011;
            15'd20440: log10_cal = 16'b0000010100110011;
            15'd20441: log10_cal = 16'b0000010100110011;
            15'd20442: log10_cal = 16'b0000010100110011;
            15'd20443: log10_cal = 16'b0000010100110011;
            15'd20444: log10_cal = 16'b0000010100110011;
            15'd20445: log10_cal = 16'b0000010100110011;
            15'd20446: log10_cal = 16'b0000010100110011;
            15'd20447: log10_cal = 16'b0000010100110011;
            15'd20448: log10_cal = 16'b0000010100110011;
            15'd20449: log10_cal = 16'b0000010100110011;
            15'd20450: log10_cal = 16'b0000010100110011;
            15'd20451: log10_cal = 16'b0000010100110011;
            15'd20452: log10_cal = 16'b0000010100110011;
            15'd20453: log10_cal = 16'b0000010100110011;
            15'd20454: log10_cal = 16'b0000010100110011;
            15'd20455: log10_cal = 16'b0000010100110011;
            15'd20456: log10_cal = 16'b0000010100110011;
            15'd20457: log10_cal = 16'b0000010100110011;
            15'd20458: log10_cal = 16'b0000010100110011;
            15'd20459: log10_cal = 16'b0000010100110011;
            15'd20460: log10_cal = 16'b0000010100110011;
            15'd20461: log10_cal = 16'b0000010100110011;
            15'd20462: log10_cal = 16'b0000010100110011;
            15'd20463: log10_cal = 16'b0000010100110011;
            15'd20464: log10_cal = 16'b0000010100110011;
            15'd20465: log10_cal = 16'b0000010100110011;
            15'd20466: log10_cal = 16'b0000010100110011;
            15'd20467: log10_cal = 16'b0000010100110011;
            15'd20468: log10_cal = 16'b0000010100110011;
            15'd20469: log10_cal = 16'b0000010100110100;
            15'd20470: log10_cal = 16'b0000010100110100;
            15'd20471: log10_cal = 16'b0000010100110100;
            15'd20472: log10_cal = 16'b0000010100110100;
            15'd20473: log10_cal = 16'b0000010100110100;
            15'd20474: log10_cal = 16'b0000010100110100;
            15'd20475: log10_cal = 16'b0000010100110100;
            15'd20476: log10_cal = 16'b0000010100110100;
            15'd20477: log10_cal = 16'b0000010100110100;
            15'd20478: log10_cal = 16'b0000010100110100;
            15'd20479: log10_cal = 16'b0000010100110100;
            15'd20480: log10_cal = 16'b0000010100110100;
            15'd20481: log10_cal = 16'b0000010100110100;
            15'd20482: log10_cal = 16'b0000010100110100;
            15'd20483: log10_cal = 16'b0000010100110100;
            15'd20484: log10_cal = 16'b0000010100110100;
            15'd20485: log10_cal = 16'b0000010100110100;
            15'd20486: log10_cal = 16'b0000010100110100;
            15'd20487: log10_cal = 16'b0000010100110100;
            15'd20488: log10_cal = 16'b0000010100110100;
            15'd20489: log10_cal = 16'b0000010100110100;
            15'd20490: log10_cal = 16'b0000010100110100;
            15'd20491: log10_cal = 16'b0000010100110100;
            15'd20492: log10_cal = 16'b0000010100110100;
            15'd20493: log10_cal = 16'b0000010100110100;
            15'd20494: log10_cal = 16'b0000010100110100;
            15'd20495: log10_cal = 16'b0000010100110100;
            15'd20496: log10_cal = 16'b0000010100110100;
            15'd20497: log10_cal = 16'b0000010100110100;
            15'd20498: log10_cal = 16'b0000010100110100;
            15'd20499: log10_cal = 16'b0000010100110100;
            15'd20500: log10_cal = 16'b0000010100110100;
            15'd20501: log10_cal = 16'b0000010100110100;
            15'd20502: log10_cal = 16'b0000010100110100;
            15'd20503: log10_cal = 16'b0000010100110100;
            15'd20504: log10_cal = 16'b0000010100110100;
            15'd20505: log10_cal = 16'b0000010100110100;
            15'd20506: log10_cal = 16'b0000010100110100;
            15'd20507: log10_cal = 16'b0000010100110100;
            15'd20508: log10_cal = 16'b0000010100110100;
            15'd20509: log10_cal = 16'b0000010100110100;
            15'd20510: log10_cal = 16'b0000010100110100;
            15'd20511: log10_cal = 16'b0000010100110100;
            15'd20512: log10_cal = 16'b0000010100110100;
            15'd20513: log10_cal = 16'b0000010100110100;
            15'd20514: log10_cal = 16'b0000010100110100;
            15'd20515: log10_cal = 16'b0000010100110101;
            15'd20516: log10_cal = 16'b0000010100110101;
            15'd20517: log10_cal = 16'b0000010100110101;
            15'd20518: log10_cal = 16'b0000010100110101;
            15'd20519: log10_cal = 16'b0000010100110101;
            15'd20520: log10_cal = 16'b0000010100110101;
            15'd20521: log10_cal = 16'b0000010100110101;
            15'd20522: log10_cal = 16'b0000010100110101;
            15'd20523: log10_cal = 16'b0000010100110101;
            15'd20524: log10_cal = 16'b0000010100110101;
            15'd20525: log10_cal = 16'b0000010100110101;
            15'd20526: log10_cal = 16'b0000010100110101;
            15'd20527: log10_cal = 16'b0000010100110101;
            15'd20528: log10_cal = 16'b0000010100110101;
            15'd20529: log10_cal = 16'b0000010100110101;
            15'd20530: log10_cal = 16'b0000010100110101;
            15'd20531: log10_cal = 16'b0000010100110101;
            15'd20532: log10_cal = 16'b0000010100110101;
            15'd20533: log10_cal = 16'b0000010100110101;
            15'd20534: log10_cal = 16'b0000010100110101;
            15'd20535: log10_cal = 16'b0000010100110101;
            15'd20536: log10_cal = 16'b0000010100110101;
            15'd20537: log10_cal = 16'b0000010100110101;
            15'd20538: log10_cal = 16'b0000010100110101;
            15'd20539: log10_cal = 16'b0000010100110101;
            15'd20540: log10_cal = 16'b0000010100110101;
            15'd20541: log10_cal = 16'b0000010100110101;
            15'd20542: log10_cal = 16'b0000010100110101;
            15'd20543: log10_cal = 16'b0000010100110101;
            15'd20544: log10_cal = 16'b0000010100110101;
            15'd20545: log10_cal = 16'b0000010100110101;
            15'd20546: log10_cal = 16'b0000010100110101;
            15'd20547: log10_cal = 16'b0000010100110101;
            15'd20548: log10_cal = 16'b0000010100110101;
            15'd20549: log10_cal = 16'b0000010100110101;
            15'd20550: log10_cal = 16'b0000010100110101;
            15'd20551: log10_cal = 16'b0000010100110101;
            15'd20552: log10_cal = 16'b0000010100110101;
            15'd20553: log10_cal = 16'b0000010100110101;
            15'd20554: log10_cal = 16'b0000010100110101;
            15'd20555: log10_cal = 16'b0000010100110101;
            15'd20556: log10_cal = 16'b0000010100110101;
            15'd20557: log10_cal = 16'b0000010100110101;
            15'd20558: log10_cal = 16'b0000010100110101;
            15'd20559: log10_cal = 16'b0000010100110101;
            15'd20560: log10_cal = 16'b0000010100110101;
            15'd20561: log10_cal = 16'b0000010100110110;
            15'd20562: log10_cal = 16'b0000010100110110;
            15'd20563: log10_cal = 16'b0000010100110110;
            15'd20564: log10_cal = 16'b0000010100110110;
            15'd20565: log10_cal = 16'b0000010100110110;
            15'd20566: log10_cal = 16'b0000010100110110;
            15'd20567: log10_cal = 16'b0000010100110110;
            15'd20568: log10_cal = 16'b0000010100110110;
            15'd20569: log10_cal = 16'b0000010100110110;
            15'd20570: log10_cal = 16'b0000010100110110;
            15'd20571: log10_cal = 16'b0000010100110110;
            15'd20572: log10_cal = 16'b0000010100110110;
            15'd20573: log10_cal = 16'b0000010100110110;
            15'd20574: log10_cal = 16'b0000010100110110;
            15'd20575: log10_cal = 16'b0000010100110110;
            15'd20576: log10_cal = 16'b0000010100110110;
            15'd20577: log10_cal = 16'b0000010100110110;
            15'd20578: log10_cal = 16'b0000010100110110;
            15'd20579: log10_cal = 16'b0000010100110110;
            15'd20580: log10_cal = 16'b0000010100110110;
            15'd20581: log10_cal = 16'b0000010100110110;
            15'd20582: log10_cal = 16'b0000010100110110;
            15'd20583: log10_cal = 16'b0000010100110110;
            15'd20584: log10_cal = 16'b0000010100110110;
            15'd20585: log10_cal = 16'b0000010100110110;
            15'd20586: log10_cal = 16'b0000010100110110;
            15'd20587: log10_cal = 16'b0000010100110110;
            15'd20588: log10_cal = 16'b0000010100110110;
            15'd20589: log10_cal = 16'b0000010100110110;
            15'd20590: log10_cal = 16'b0000010100110110;
            15'd20591: log10_cal = 16'b0000010100110110;
            15'd20592: log10_cal = 16'b0000010100110110;
            15'd20593: log10_cal = 16'b0000010100110110;
            15'd20594: log10_cal = 16'b0000010100110110;
            15'd20595: log10_cal = 16'b0000010100110110;
            15'd20596: log10_cal = 16'b0000010100110110;
            15'd20597: log10_cal = 16'b0000010100110110;
            15'd20598: log10_cal = 16'b0000010100110110;
            15'd20599: log10_cal = 16'b0000010100110110;
            15'd20600: log10_cal = 16'b0000010100110110;
            15'd20601: log10_cal = 16'b0000010100110110;
            15'd20602: log10_cal = 16'b0000010100110110;
            15'd20603: log10_cal = 16'b0000010100110110;
            15'd20604: log10_cal = 16'b0000010100110110;
            15'd20605: log10_cal = 16'b0000010100110110;
            15'd20606: log10_cal = 16'b0000010100110110;
            15'd20607: log10_cal = 16'b0000010100110111;
            15'd20608: log10_cal = 16'b0000010100110111;
            15'd20609: log10_cal = 16'b0000010100110111;
            15'd20610: log10_cal = 16'b0000010100110111;
            15'd20611: log10_cal = 16'b0000010100110111;
            15'd20612: log10_cal = 16'b0000010100110111;
            15'd20613: log10_cal = 16'b0000010100110111;
            15'd20614: log10_cal = 16'b0000010100110111;
            15'd20615: log10_cal = 16'b0000010100110111;
            15'd20616: log10_cal = 16'b0000010100110111;
            15'd20617: log10_cal = 16'b0000010100110111;
            15'd20618: log10_cal = 16'b0000010100110111;
            15'd20619: log10_cal = 16'b0000010100110111;
            15'd20620: log10_cal = 16'b0000010100110111;
            15'd20621: log10_cal = 16'b0000010100110111;
            15'd20622: log10_cal = 16'b0000010100110111;
            15'd20623: log10_cal = 16'b0000010100110111;
            15'd20624: log10_cal = 16'b0000010100110111;
            15'd20625: log10_cal = 16'b0000010100110111;
            15'd20626: log10_cal = 16'b0000010100110111;
            15'd20627: log10_cal = 16'b0000010100110111;
            15'd20628: log10_cal = 16'b0000010100110111;
            15'd20629: log10_cal = 16'b0000010100110111;
            15'd20630: log10_cal = 16'b0000010100110111;
            15'd20631: log10_cal = 16'b0000010100110111;
            15'd20632: log10_cal = 16'b0000010100110111;
            15'd20633: log10_cal = 16'b0000010100110111;
            15'd20634: log10_cal = 16'b0000010100110111;
            15'd20635: log10_cal = 16'b0000010100110111;
            15'd20636: log10_cal = 16'b0000010100110111;
            15'd20637: log10_cal = 16'b0000010100110111;
            15'd20638: log10_cal = 16'b0000010100110111;
            15'd20639: log10_cal = 16'b0000010100110111;
            15'd20640: log10_cal = 16'b0000010100110111;
            15'd20641: log10_cal = 16'b0000010100110111;
            15'd20642: log10_cal = 16'b0000010100110111;
            15'd20643: log10_cal = 16'b0000010100110111;
            15'd20644: log10_cal = 16'b0000010100110111;
            15'd20645: log10_cal = 16'b0000010100110111;
            15'd20646: log10_cal = 16'b0000010100110111;
            15'd20647: log10_cal = 16'b0000010100110111;
            15'd20648: log10_cal = 16'b0000010100110111;
            15'd20649: log10_cal = 16'b0000010100110111;
            15'd20650: log10_cal = 16'b0000010100110111;
            15'd20651: log10_cal = 16'b0000010100110111;
            15'd20652: log10_cal = 16'b0000010100110111;
            15'd20653: log10_cal = 16'b0000010100110111;
            15'd20654: log10_cal = 16'b0000010100111000;
            15'd20655: log10_cal = 16'b0000010100111000;
            15'd20656: log10_cal = 16'b0000010100111000;
            15'd20657: log10_cal = 16'b0000010100111000;
            15'd20658: log10_cal = 16'b0000010100111000;
            15'd20659: log10_cal = 16'b0000010100111000;
            15'd20660: log10_cal = 16'b0000010100111000;
            15'd20661: log10_cal = 16'b0000010100111000;
            15'd20662: log10_cal = 16'b0000010100111000;
            15'd20663: log10_cal = 16'b0000010100111000;
            15'd20664: log10_cal = 16'b0000010100111000;
            15'd20665: log10_cal = 16'b0000010100111000;
            15'd20666: log10_cal = 16'b0000010100111000;
            15'd20667: log10_cal = 16'b0000010100111000;
            15'd20668: log10_cal = 16'b0000010100111000;
            15'd20669: log10_cal = 16'b0000010100111000;
            15'd20670: log10_cal = 16'b0000010100111000;
            15'd20671: log10_cal = 16'b0000010100111000;
            15'd20672: log10_cal = 16'b0000010100111000;
            15'd20673: log10_cal = 16'b0000010100111000;
            15'd20674: log10_cal = 16'b0000010100111000;
            15'd20675: log10_cal = 16'b0000010100111000;
            15'd20676: log10_cal = 16'b0000010100111000;
            15'd20677: log10_cal = 16'b0000010100111000;
            15'd20678: log10_cal = 16'b0000010100111000;
            15'd20679: log10_cal = 16'b0000010100111000;
            15'd20680: log10_cal = 16'b0000010100111000;
            15'd20681: log10_cal = 16'b0000010100111000;
            15'd20682: log10_cal = 16'b0000010100111000;
            15'd20683: log10_cal = 16'b0000010100111000;
            15'd20684: log10_cal = 16'b0000010100111000;
            15'd20685: log10_cal = 16'b0000010100111000;
            15'd20686: log10_cal = 16'b0000010100111000;
            15'd20687: log10_cal = 16'b0000010100111000;
            15'd20688: log10_cal = 16'b0000010100111000;
            15'd20689: log10_cal = 16'b0000010100111000;
            15'd20690: log10_cal = 16'b0000010100111000;
            15'd20691: log10_cal = 16'b0000010100111000;
            15'd20692: log10_cal = 16'b0000010100111000;
            15'd20693: log10_cal = 16'b0000010100111000;
            15'd20694: log10_cal = 16'b0000010100111000;
            15'd20695: log10_cal = 16'b0000010100111000;
            15'd20696: log10_cal = 16'b0000010100111000;
            15'd20697: log10_cal = 16'b0000010100111000;
            15'd20698: log10_cal = 16'b0000010100111000;
            15'd20699: log10_cal = 16'b0000010100111000;
            15'd20700: log10_cal = 16'b0000010100111001;
            15'd20701: log10_cal = 16'b0000010100111001;
            15'd20702: log10_cal = 16'b0000010100111001;
            15'd20703: log10_cal = 16'b0000010100111001;
            15'd20704: log10_cal = 16'b0000010100111001;
            15'd20705: log10_cal = 16'b0000010100111001;
            15'd20706: log10_cal = 16'b0000010100111001;
            15'd20707: log10_cal = 16'b0000010100111001;
            15'd20708: log10_cal = 16'b0000010100111001;
            15'd20709: log10_cal = 16'b0000010100111001;
            15'd20710: log10_cal = 16'b0000010100111001;
            15'd20711: log10_cal = 16'b0000010100111001;
            15'd20712: log10_cal = 16'b0000010100111001;
            15'd20713: log10_cal = 16'b0000010100111001;
            15'd20714: log10_cal = 16'b0000010100111001;
            15'd20715: log10_cal = 16'b0000010100111001;
            15'd20716: log10_cal = 16'b0000010100111001;
            15'd20717: log10_cal = 16'b0000010100111001;
            15'd20718: log10_cal = 16'b0000010100111001;
            15'd20719: log10_cal = 16'b0000010100111001;
            15'd20720: log10_cal = 16'b0000010100111001;
            15'd20721: log10_cal = 16'b0000010100111001;
            15'd20722: log10_cal = 16'b0000010100111001;
            15'd20723: log10_cal = 16'b0000010100111001;
            15'd20724: log10_cal = 16'b0000010100111001;
            15'd20725: log10_cal = 16'b0000010100111001;
            15'd20726: log10_cal = 16'b0000010100111001;
            15'd20727: log10_cal = 16'b0000010100111001;
            15'd20728: log10_cal = 16'b0000010100111001;
            15'd20729: log10_cal = 16'b0000010100111001;
            15'd20730: log10_cal = 16'b0000010100111001;
            15'd20731: log10_cal = 16'b0000010100111001;
            15'd20732: log10_cal = 16'b0000010100111001;
            15'd20733: log10_cal = 16'b0000010100111001;
            15'd20734: log10_cal = 16'b0000010100111001;
            15'd20735: log10_cal = 16'b0000010100111001;
            15'd20736: log10_cal = 16'b0000010100111001;
            15'd20737: log10_cal = 16'b0000010100111001;
            15'd20738: log10_cal = 16'b0000010100111001;
            15'd20739: log10_cal = 16'b0000010100111001;
            15'd20740: log10_cal = 16'b0000010100111001;
            15'd20741: log10_cal = 16'b0000010100111001;
            15'd20742: log10_cal = 16'b0000010100111001;
            15'd20743: log10_cal = 16'b0000010100111001;
            15'd20744: log10_cal = 16'b0000010100111001;
            15'd20745: log10_cal = 16'b0000010100111001;
            15'd20746: log10_cal = 16'b0000010100111001;
            15'd20747: log10_cal = 16'b0000010100111010;
            15'd20748: log10_cal = 16'b0000010100111010;
            15'd20749: log10_cal = 16'b0000010100111010;
            15'd20750: log10_cal = 16'b0000010100111010;
            15'd20751: log10_cal = 16'b0000010100111010;
            15'd20752: log10_cal = 16'b0000010100111010;
            15'd20753: log10_cal = 16'b0000010100111010;
            15'd20754: log10_cal = 16'b0000010100111010;
            15'd20755: log10_cal = 16'b0000010100111010;
            15'd20756: log10_cal = 16'b0000010100111010;
            15'd20757: log10_cal = 16'b0000010100111010;
            15'd20758: log10_cal = 16'b0000010100111010;
            15'd20759: log10_cal = 16'b0000010100111010;
            15'd20760: log10_cal = 16'b0000010100111010;
            15'd20761: log10_cal = 16'b0000010100111010;
            15'd20762: log10_cal = 16'b0000010100111010;
            15'd20763: log10_cal = 16'b0000010100111010;
            15'd20764: log10_cal = 16'b0000010100111010;
            15'd20765: log10_cal = 16'b0000010100111010;
            15'd20766: log10_cal = 16'b0000010100111010;
            15'd20767: log10_cal = 16'b0000010100111010;
            15'd20768: log10_cal = 16'b0000010100111010;
            15'd20769: log10_cal = 16'b0000010100111010;
            15'd20770: log10_cal = 16'b0000010100111010;
            15'd20771: log10_cal = 16'b0000010100111010;
            15'd20772: log10_cal = 16'b0000010100111010;
            15'd20773: log10_cal = 16'b0000010100111010;
            15'd20774: log10_cal = 16'b0000010100111010;
            15'd20775: log10_cal = 16'b0000010100111010;
            15'd20776: log10_cal = 16'b0000010100111010;
            15'd20777: log10_cal = 16'b0000010100111010;
            15'd20778: log10_cal = 16'b0000010100111010;
            15'd20779: log10_cal = 16'b0000010100111010;
            15'd20780: log10_cal = 16'b0000010100111010;
            15'd20781: log10_cal = 16'b0000010100111010;
            15'd20782: log10_cal = 16'b0000010100111010;
            15'd20783: log10_cal = 16'b0000010100111010;
            15'd20784: log10_cal = 16'b0000010100111010;
            15'd20785: log10_cal = 16'b0000010100111010;
            15'd20786: log10_cal = 16'b0000010100111010;
            15'd20787: log10_cal = 16'b0000010100111010;
            15'd20788: log10_cal = 16'b0000010100111010;
            15'd20789: log10_cal = 16'b0000010100111010;
            15'd20790: log10_cal = 16'b0000010100111010;
            15'd20791: log10_cal = 16'b0000010100111010;
            15'd20792: log10_cal = 16'b0000010100111010;
            15'd20793: log10_cal = 16'b0000010100111011;
            15'd20794: log10_cal = 16'b0000010100111011;
            15'd20795: log10_cal = 16'b0000010100111011;
            15'd20796: log10_cal = 16'b0000010100111011;
            15'd20797: log10_cal = 16'b0000010100111011;
            15'd20798: log10_cal = 16'b0000010100111011;
            15'd20799: log10_cal = 16'b0000010100111011;
            15'd20800: log10_cal = 16'b0000010100111011;
            15'd20801: log10_cal = 16'b0000010100111011;
            15'd20802: log10_cal = 16'b0000010100111011;
            15'd20803: log10_cal = 16'b0000010100111011;
            15'd20804: log10_cal = 16'b0000010100111011;
            15'd20805: log10_cal = 16'b0000010100111011;
            15'd20806: log10_cal = 16'b0000010100111011;
            15'd20807: log10_cal = 16'b0000010100111011;
            15'd20808: log10_cal = 16'b0000010100111011;
            15'd20809: log10_cal = 16'b0000010100111011;
            15'd20810: log10_cal = 16'b0000010100111011;
            15'd20811: log10_cal = 16'b0000010100111011;
            15'd20812: log10_cal = 16'b0000010100111011;
            15'd20813: log10_cal = 16'b0000010100111011;
            15'd20814: log10_cal = 16'b0000010100111011;
            15'd20815: log10_cal = 16'b0000010100111011;
            15'd20816: log10_cal = 16'b0000010100111011;
            15'd20817: log10_cal = 16'b0000010100111011;
            15'd20818: log10_cal = 16'b0000010100111011;
            15'd20819: log10_cal = 16'b0000010100111011;
            15'd20820: log10_cal = 16'b0000010100111011;
            15'd20821: log10_cal = 16'b0000010100111011;
            15'd20822: log10_cal = 16'b0000010100111011;
            15'd20823: log10_cal = 16'b0000010100111011;
            15'd20824: log10_cal = 16'b0000010100111011;
            15'd20825: log10_cal = 16'b0000010100111011;
            15'd20826: log10_cal = 16'b0000010100111011;
            15'd20827: log10_cal = 16'b0000010100111011;
            15'd20828: log10_cal = 16'b0000010100111011;
            15'd20829: log10_cal = 16'b0000010100111011;
            15'd20830: log10_cal = 16'b0000010100111011;
            15'd20831: log10_cal = 16'b0000010100111011;
            15'd20832: log10_cal = 16'b0000010100111011;
            15'd20833: log10_cal = 16'b0000010100111011;
            15'd20834: log10_cal = 16'b0000010100111011;
            15'd20835: log10_cal = 16'b0000010100111011;
            15'd20836: log10_cal = 16'b0000010100111011;
            15'd20837: log10_cal = 16'b0000010100111011;
            15'd20838: log10_cal = 16'b0000010100111011;
            15'd20839: log10_cal = 16'b0000010100111011;
            15'd20840: log10_cal = 16'b0000010100111100;
            15'd20841: log10_cal = 16'b0000010100111100;
            15'd20842: log10_cal = 16'b0000010100111100;
            15'd20843: log10_cal = 16'b0000010100111100;
            15'd20844: log10_cal = 16'b0000010100111100;
            15'd20845: log10_cal = 16'b0000010100111100;
            15'd20846: log10_cal = 16'b0000010100111100;
            15'd20847: log10_cal = 16'b0000010100111100;
            15'd20848: log10_cal = 16'b0000010100111100;
            15'd20849: log10_cal = 16'b0000010100111100;
            15'd20850: log10_cal = 16'b0000010100111100;
            15'd20851: log10_cal = 16'b0000010100111100;
            15'd20852: log10_cal = 16'b0000010100111100;
            15'd20853: log10_cal = 16'b0000010100111100;
            15'd20854: log10_cal = 16'b0000010100111100;
            15'd20855: log10_cal = 16'b0000010100111100;
            15'd20856: log10_cal = 16'b0000010100111100;
            15'd20857: log10_cal = 16'b0000010100111100;
            15'd20858: log10_cal = 16'b0000010100111100;
            15'd20859: log10_cal = 16'b0000010100111100;
            15'd20860: log10_cal = 16'b0000010100111100;
            15'd20861: log10_cal = 16'b0000010100111100;
            15'd20862: log10_cal = 16'b0000010100111100;
            15'd20863: log10_cal = 16'b0000010100111100;
            15'd20864: log10_cal = 16'b0000010100111100;
            15'd20865: log10_cal = 16'b0000010100111100;
            15'd20866: log10_cal = 16'b0000010100111100;
            15'd20867: log10_cal = 16'b0000010100111100;
            15'd20868: log10_cal = 16'b0000010100111100;
            15'd20869: log10_cal = 16'b0000010100111100;
            15'd20870: log10_cal = 16'b0000010100111100;
            15'd20871: log10_cal = 16'b0000010100111100;
            15'd20872: log10_cal = 16'b0000010100111100;
            15'd20873: log10_cal = 16'b0000010100111100;
            15'd20874: log10_cal = 16'b0000010100111100;
            15'd20875: log10_cal = 16'b0000010100111100;
            15'd20876: log10_cal = 16'b0000010100111100;
            15'd20877: log10_cal = 16'b0000010100111100;
            15'd20878: log10_cal = 16'b0000010100111100;
            15'd20879: log10_cal = 16'b0000010100111100;
            15'd20880: log10_cal = 16'b0000010100111100;
            15'd20881: log10_cal = 16'b0000010100111100;
            15'd20882: log10_cal = 16'b0000010100111100;
            15'd20883: log10_cal = 16'b0000010100111100;
            15'd20884: log10_cal = 16'b0000010100111100;
            15'd20885: log10_cal = 16'b0000010100111100;
            15'd20886: log10_cal = 16'b0000010100111100;
            15'd20887: log10_cal = 16'b0000010100111101;
            15'd20888: log10_cal = 16'b0000010100111101;
            15'd20889: log10_cal = 16'b0000010100111101;
            15'd20890: log10_cal = 16'b0000010100111101;
            15'd20891: log10_cal = 16'b0000010100111101;
            15'd20892: log10_cal = 16'b0000010100111101;
            15'd20893: log10_cal = 16'b0000010100111101;
            15'd20894: log10_cal = 16'b0000010100111101;
            15'd20895: log10_cal = 16'b0000010100111101;
            15'd20896: log10_cal = 16'b0000010100111101;
            15'd20897: log10_cal = 16'b0000010100111101;
            15'd20898: log10_cal = 16'b0000010100111101;
            15'd20899: log10_cal = 16'b0000010100111101;
            15'd20900: log10_cal = 16'b0000010100111101;
            15'd20901: log10_cal = 16'b0000010100111101;
            15'd20902: log10_cal = 16'b0000010100111101;
            15'd20903: log10_cal = 16'b0000010100111101;
            15'd20904: log10_cal = 16'b0000010100111101;
            15'd20905: log10_cal = 16'b0000010100111101;
            15'd20906: log10_cal = 16'b0000010100111101;
            15'd20907: log10_cal = 16'b0000010100111101;
            15'd20908: log10_cal = 16'b0000010100111101;
            15'd20909: log10_cal = 16'b0000010100111101;
            15'd20910: log10_cal = 16'b0000010100111101;
            15'd20911: log10_cal = 16'b0000010100111101;
            15'd20912: log10_cal = 16'b0000010100111101;
            15'd20913: log10_cal = 16'b0000010100111101;
            15'd20914: log10_cal = 16'b0000010100111101;
            15'd20915: log10_cal = 16'b0000010100111101;
            15'd20916: log10_cal = 16'b0000010100111101;
            15'd20917: log10_cal = 16'b0000010100111101;
            15'd20918: log10_cal = 16'b0000010100111101;
            15'd20919: log10_cal = 16'b0000010100111101;
            15'd20920: log10_cal = 16'b0000010100111101;
            15'd20921: log10_cal = 16'b0000010100111101;
            15'd20922: log10_cal = 16'b0000010100111101;
            15'd20923: log10_cal = 16'b0000010100111101;
            15'd20924: log10_cal = 16'b0000010100111101;
            15'd20925: log10_cal = 16'b0000010100111101;
            15'd20926: log10_cal = 16'b0000010100111101;
            15'd20927: log10_cal = 16'b0000010100111101;
            15'd20928: log10_cal = 16'b0000010100111101;
            15'd20929: log10_cal = 16'b0000010100111101;
            15'd20930: log10_cal = 16'b0000010100111101;
            15'd20931: log10_cal = 16'b0000010100111101;
            15'd20932: log10_cal = 16'b0000010100111101;
            15'd20933: log10_cal = 16'b0000010100111101;
            15'd20934: log10_cal = 16'b0000010100111110;
            15'd20935: log10_cal = 16'b0000010100111110;
            15'd20936: log10_cal = 16'b0000010100111110;
            15'd20937: log10_cal = 16'b0000010100111110;
            15'd20938: log10_cal = 16'b0000010100111110;
            15'd20939: log10_cal = 16'b0000010100111110;
            15'd20940: log10_cal = 16'b0000010100111110;
            15'd20941: log10_cal = 16'b0000010100111110;
            15'd20942: log10_cal = 16'b0000010100111110;
            15'd20943: log10_cal = 16'b0000010100111110;
            15'd20944: log10_cal = 16'b0000010100111110;
            15'd20945: log10_cal = 16'b0000010100111110;
            15'd20946: log10_cal = 16'b0000010100111110;
            15'd20947: log10_cal = 16'b0000010100111110;
            15'd20948: log10_cal = 16'b0000010100111110;
            15'd20949: log10_cal = 16'b0000010100111110;
            15'd20950: log10_cal = 16'b0000010100111110;
            15'd20951: log10_cal = 16'b0000010100111110;
            15'd20952: log10_cal = 16'b0000010100111110;
            15'd20953: log10_cal = 16'b0000010100111110;
            15'd20954: log10_cal = 16'b0000010100111110;
            15'd20955: log10_cal = 16'b0000010100111110;
            15'd20956: log10_cal = 16'b0000010100111110;
            15'd20957: log10_cal = 16'b0000010100111110;
            15'd20958: log10_cal = 16'b0000010100111110;
            15'd20959: log10_cal = 16'b0000010100111110;
            15'd20960: log10_cal = 16'b0000010100111110;
            15'd20961: log10_cal = 16'b0000010100111110;
            15'd20962: log10_cal = 16'b0000010100111110;
            15'd20963: log10_cal = 16'b0000010100111110;
            15'd20964: log10_cal = 16'b0000010100111110;
            15'd20965: log10_cal = 16'b0000010100111110;
            15'd20966: log10_cal = 16'b0000010100111110;
            15'd20967: log10_cal = 16'b0000010100111110;
            15'd20968: log10_cal = 16'b0000010100111110;
            15'd20969: log10_cal = 16'b0000010100111110;
            15'd20970: log10_cal = 16'b0000010100111110;
            15'd20971: log10_cal = 16'b0000010100111110;
            15'd20972: log10_cal = 16'b0000010100111110;
            15'd20973: log10_cal = 16'b0000010100111110;
            15'd20974: log10_cal = 16'b0000010100111110;
            15'd20975: log10_cal = 16'b0000010100111110;
            15'd20976: log10_cal = 16'b0000010100111110;
            15'd20977: log10_cal = 16'b0000010100111110;
            15'd20978: log10_cal = 16'b0000010100111110;
            15'd20979: log10_cal = 16'b0000010100111110;
            15'd20980: log10_cal = 16'b0000010100111110;
            15'd20981: log10_cal = 16'b0000010100111111;
            15'd20982: log10_cal = 16'b0000010100111111;
            15'd20983: log10_cal = 16'b0000010100111111;
            15'd20984: log10_cal = 16'b0000010100111111;
            15'd20985: log10_cal = 16'b0000010100111111;
            15'd20986: log10_cal = 16'b0000010100111111;
            15'd20987: log10_cal = 16'b0000010100111111;
            15'd20988: log10_cal = 16'b0000010100111111;
            15'd20989: log10_cal = 16'b0000010100111111;
            15'd20990: log10_cal = 16'b0000010100111111;
            15'd20991: log10_cal = 16'b0000010100111111;
            15'd20992: log10_cal = 16'b0000010100111111;
            15'd20993: log10_cal = 16'b0000010100111111;
            15'd20994: log10_cal = 16'b0000010100111111;
            15'd20995: log10_cal = 16'b0000010100111111;
            15'd20996: log10_cal = 16'b0000010100111111;
            15'd20997: log10_cal = 16'b0000010100111111;
            15'd20998: log10_cal = 16'b0000010100111111;
            15'd20999: log10_cal = 16'b0000010100111111;
            15'd21000: log10_cal = 16'b0000010100111111;
            15'd21001: log10_cal = 16'b0000010100111111;
            15'd21002: log10_cal = 16'b0000010100111111;
            15'd21003: log10_cal = 16'b0000010100111111;
            15'd21004: log10_cal = 16'b0000010100111111;
            15'd21005: log10_cal = 16'b0000010100111111;
            15'd21006: log10_cal = 16'b0000010100111111;
            15'd21007: log10_cal = 16'b0000010100111111;
            15'd21008: log10_cal = 16'b0000010100111111;
            15'd21009: log10_cal = 16'b0000010100111111;
            15'd21010: log10_cal = 16'b0000010100111111;
            15'd21011: log10_cal = 16'b0000010100111111;
            15'd21012: log10_cal = 16'b0000010100111111;
            15'd21013: log10_cal = 16'b0000010100111111;
            15'd21014: log10_cal = 16'b0000010100111111;
            15'd21015: log10_cal = 16'b0000010100111111;
            15'd21016: log10_cal = 16'b0000010100111111;
            15'd21017: log10_cal = 16'b0000010100111111;
            15'd21018: log10_cal = 16'b0000010100111111;
            15'd21019: log10_cal = 16'b0000010100111111;
            15'd21020: log10_cal = 16'b0000010100111111;
            15'd21021: log10_cal = 16'b0000010100111111;
            15'd21022: log10_cal = 16'b0000010100111111;
            15'd21023: log10_cal = 16'b0000010100111111;
            15'd21024: log10_cal = 16'b0000010100111111;
            15'd21025: log10_cal = 16'b0000010100111111;
            15'd21026: log10_cal = 16'b0000010100111111;
            15'd21027: log10_cal = 16'b0000010100111111;
            15'd21028: log10_cal = 16'b0000010100111111;
            15'd21029: log10_cal = 16'b0000010101000000;
            15'd21030: log10_cal = 16'b0000010101000000;
            15'd21031: log10_cal = 16'b0000010101000000;
            15'd21032: log10_cal = 16'b0000010101000000;
            15'd21033: log10_cal = 16'b0000010101000000;
            15'd21034: log10_cal = 16'b0000010101000000;
            15'd21035: log10_cal = 16'b0000010101000000;
            15'd21036: log10_cal = 16'b0000010101000000;
            15'd21037: log10_cal = 16'b0000010101000000;
            15'd21038: log10_cal = 16'b0000010101000000;
            15'd21039: log10_cal = 16'b0000010101000000;
            15'd21040: log10_cal = 16'b0000010101000000;
            15'd21041: log10_cal = 16'b0000010101000000;
            15'd21042: log10_cal = 16'b0000010101000000;
            15'd21043: log10_cal = 16'b0000010101000000;
            15'd21044: log10_cal = 16'b0000010101000000;
            15'd21045: log10_cal = 16'b0000010101000000;
            15'd21046: log10_cal = 16'b0000010101000000;
            15'd21047: log10_cal = 16'b0000010101000000;
            15'd21048: log10_cal = 16'b0000010101000000;
            15'd21049: log10_cal = 16'b0000010101000000;
            15'd21050: log10_cal = 16'b0000010101000000;
            15'd21051: log10_cal = 16'b0000010101000000;
            15'd21052: log10_cal = 16'b0000010101000000;
            15'd21053: log10_cal = 16'b0000010101000000;
            15'd21054: log10_cal = 16'b0000010101000000;
            15'd21055: log10_cal = 16'b0000010101000000;
            15'd21056: log10_cal = 16'b0000010101000000;
            15'd21057: log10_cal = 16'b0000010101000000;
            15'd21058: log10_cal = 16'b0000010101000000;
            15'd21059: log10_cal = 16'b0000010101000000;
            15'd21060: log10_cal = 16'b0000010101000000;
            15'd21061: log10_cal = 16'b0000010101000000;
            15'd21062: log10_cal = 16'b0000010101000000;
            15'd21063: log10_cal = 16'b0000010101000000;
            15'd21064: log10_cal = 16'b0000010101000000;
            15'd21065: log10_cal = 16'b0000010101000000;
            15'd21066: log10_cal = 16'b0000010101000000;
            15'd21067: log10_cal = 16'b0000010101000000;
            15'd21068: log10_cal = 16'b0000010101000000;
            15'd21069: log10_cal = 16'b0000010101000000;
            15'd21070: log10_cal = 16'b0000010101000000;
            15'd21071: log10_cal = 16'b0000010101000000;
            15'd21072: log10_cal = 16'b0000010101000000;
            15'd21073: log10_cal = 16'b0000010101000000;
            15'd21074: log10_cal = 16'b0000010101000000;
            15'd21075: log10_cal = 16'b0000010101000000;
            15'd21076: log10_cal = 16'b0000010101000001;
            15'd21077: log10_cal = 16'b0000010101000001;
            15'd21078: log10_cal = 16'b0000010101000001;
            15'd21079: log10_cal = 16'b0000010101000001;
            15'd21080: log10_cal = 16'b0000010101000001;
            15'd21081: log10_cal = 16'b0000010101000001;
            15'd21082: log10_cal = 16'b0000010101000001;
            15'd21083: log10_cal = 16'b0000010101000001;
            15'd21084: log10_cal = 16'b0000010101000001;
            15'd21085: log10_cal = 16'b0000010101000001;
            15'd21086: log10_cal = 16'b0000010101000001;
            15'd21087: log10_cal = 16'b0000010101000001;
            15'd21088: log10_cal = 16'b0000010101000001;
            15'd21089: log10_cal = 16'b0000010101000001;
            15'd21090: log10_cal = 16'b0000010101000001;
            15'd21091: log10_cal = 16'b0000010101000001;
            15'd21092: log10_cal = 16'b0000010101000001;
            15'd21093: log10_cal = 16'b0000010101000001;
            15'd21094: log10_cal = 16'b0000010101000001;
            15'd21095: log10_cal = 16'b0000010101000001;
            15'd21096: log10_cal = 16'b0000010101000001;
            15'd21097: log10_cal = 16'b0000010101000001;
            15'd21098: log10_cal = 16'b0000010101000001;
            15'd21099: log10_cal = 16'b0000010101000001;
            15'd21100: log10_cal = 16'b0000010101000001;
            15'd21101: log10_cal = 16'b0000010101000001;
            15'd21102: log10_cal = 16'b0000010101000001;
            15'd21103: log10_cal = 16'b0000010101000001;
            15'd21104: log10_cal = 16'b0000010101000001;
            15'd21105: log10_cal = 16'b0000010101000001;
            15'd21106: log10_cal = 16'b0000010101000001;
            15'd21107: log10_cal = 16'b0000010101000001;
            15'd21108: log10_cal = 16'b0000010101000001;
            15'd21109: log10_cal = 16'b0000010101000001;
            15'd21110: log10_cal = 16'b0000010101000001;
            15'd21111: log10_cal = 16'b0000010101000001;
            15'd21112: log10_cal = 16'b0000010101000001;
            15'd21113: log10_cal = 16'b0000010101000001;
            15'd21114: log10_cal = 16'b0000010101000001;
            15'd21115: log10_cal = 16'b0000010101000001;
            15'd21116: log10_cal = 16'b0000010101000001;
            15'd21117: log10_cal = 16'b0000010101000001;
            15'd21118: log10_cal = 16'b0000010101000001;
            15'd21119: log10_cal = 16'b0000010101000001;
            15'd21120: log10_cal = 16'b0000010101000001;
            15'd21121: log10_cal = 16'b0000010101000001;
            15'd21122: log10_cal = 16'b0000010101000001;
            15'd21123: log10_cal = 16'b0000010101000010;
            15'd21124: log10_cal = 16'b0000010101000010;
            15'd21125: log10_cal = 16'b0000010101000010;
            15'd21126: log10_cal = 16'b0000010101000010;
            15'd21127: log10_cal = 16'b0000010101000010;
            15'd21128: log10_cal = 16'b0000010101000010;
            15'd21129: log10_cal = 16'b0000010101000010;
            15'd21130: log10_cal = 16'b0000010101000010;
            15'd21131: log10_cal = 16'b0000010101000010;
            15'd21132: log10_cal = 16'b0000010101000010;
            15'd21133: log10_cal = 16'b0000010101000010;
            15'd21134: log10_cal = 16'b0000010101000010;
            15'd21135: log10_cal = 16'b0000010101000010;
            15'd21136: log10_cal = 16'b0000010101000010;
            15'd21137: log10_cal = 16'b0000010101000010;
            15'd21138: log10_cal = 16'b0000010101000010;
            15'd21139: log10_cal = 16'b0000010101000010;
            15'd21140: log10_cal = 16'b0000010101000010;
            15'd21141: log10_cal = 16'b0000010101000010;
            15'd21142: log10_cal = 16'b0000010101000010;
            15'd21143: log10_cal = 16'b0000010101000010;
            15'd21144: log10_cal = 16'b0000010101000010;
            15'd21145: log10_cal = 16'b0000010101000010;
            15'd21146: log10_cal = 16'b0000010101000010;
            15'd21147: log10_cal = 16'b0000010101000010;
            15'd21148: log10_cal = 16'b0000010101000010;
            15'd21149: log10_cal = 16'b0000010101000010;
            15'd21150: log10_cal = 16'b0000010101000010;
            15'd21151: log10_cal = 16'b0000010101000010;
            15'd21152: log10_cal = 16'b0000010101000010;
            15'd21153: log10_cal = 16'b0000010101000010;
            15'd21154: log10_cal = 16'b0000010101000010;
            15'd21155: log10_cal = 16'b0000010101000010;
            15'd21156: log10_cal = 16'b0000010101000010;
            15'd21157: log10_cal = 16'b0000010101000010;
            15'd21158: log10_cal = 16'b0000010101000010;
            15'd21159: log10_cal = 16'b0000010101000010;
            15'd21160: log10_cal = 16'b0000010101000010;
            15'd21161: log10_cal = 16'b0000010101000010;
            15'd21162: log10_cal = 16'b0000010101000010;
            15'd21163: log10_cal = 16'b0000010101000010;
            15'd21164: log10_cal = 16'b0000010101000010;
            15'd21165: log10_cal = 16'b0000010101000010;
            15'd21166: log10_cal = 16'b0000010101000010;
            15'd21167: log10_cal = 16'b0000010101000010;
            15'd21168: log10_cal = 16'b0000010101000010;
            15'd21169: log10_cal = 16'b0000010101000010;
            15'd21170: log10_cal = 16'b0000010101000010;
            15'd21171: log10_cal = 16'b0000010101000011;
            15'd21172: log10_cal = 16'b0000010101000011;
            15'd21173: log10_cal = 16'b0000010101000011;
            15'd21174: log10_cal = 16'b0000010101000011;
            15'd21175: log10_cal = 16'b0000010101000011;
            15'd21176: log10_cal = 16'b0000010101000011;
            15'd21177: log10_cal = 16'b0000010101000011;
            15'd21178: log10_cal = 16'b0000010101000011;
            15'd21179: log10_cal = 16'b0000010101000011;
            15'd21180: log10_cal = 16'b0000010101000011;
            15'd21181: log10_cal = 16'b0000010101000011;
            15'd21182: log10_cal = 16'b0000010101000011;
            15'd21183: log10_cal = 16'b0000010101000011;
            15'd21184: log10_cal = 16'b0000010101000011;
            15'd21185: log10_cal = 16'b0000010101000011;
            15'd21186: log10_cal = 16'b0000010101000011;
            15'd21187: log10_cal = 16'b0000010101000011;
            15'd21188: log10_cal = 16'b0000010101000011;
            15'd21189: log10_cal = 16'b0000010101000011;
            15'd21190: log10_cal = 16'b0000010101000011;
            15'd21191: log10_cal = 16'b0000010101000011;
            15'd21192: log10_cal = 16'b0000010101000011;
            15'd21193: log10_cal = 16'b0000010101000011;
            15'd21194: log10_cal = 16'b0000010101000011;
            15'd21195: log10_cal = 16'b0000010101000011;
            15'd21196: log10_cal = 16'b0000010101000011;
            15'd21197: log10_cal = 16'b0000010101000011;
            15'd21198: log10_cal = 16'b0000010101000011;
            15'd21199: log10_cal = 16'b0000010101000011;
            15'd21200: log10_cal = 16'b0000010101000011;
            15'd21201: log10_cal = 16'b0000010101000011;
            15'd21202: log10_cal = 16'b0000010101000011;
            15'd21203: log10_cal = 16'b0000010101000011;
            15'd21204: log10_cal = 16'b0000010101000011;
            15'd21205: log10_cal = 16'b0000010101000011;
            15'd21206: log10_cal = 16'b0000010101000011;
            15'd21207: log10_cal = 16'b0000010101000011;
            15'd21208: log10_cal = 16'b0000010101000011;
            15'd21209: log10_cal = 16'b0000010101000011;
            15'd21210: log10_cal = 16'b0000010101000011;
            15'd21211: log10_cal = 16'b0000010101000011;
            15'd21212: log10_cal = 16'b0000010101000011;
            15'd21213: log10_cal = 16'b0000010101000011;
            15'd21214: log10_cal = 16'b0000010101000011;
            15'd21215: log10_cal = 16'b0000010101000011;
            15'd21216: log10_cal = 16'b0000010101000011;
            15'd21217: log10_cal = 16'b0000010101000011;
            15'd21218: log10_cal = 16'b0000010101000011;
            15'd21219: log10_cal = 16'b0000010101000100;
            15'd21220: log10_cal = 16'b0000010101000100;
            15'd21221: log10_cal = 16'b0000010101000100;
            15'd21222: log10_cal = 16'b0000010101000100;
            15'd21223: log10_cal = 16'b0000010101000100;
            15'd21224: log10_cal = 16'b0000010101000100;
            15'd21225: log10_cal = 16'b0000010101000100;
            15'd21226: log10_cal = 16'b0000010101000100;
            15'd21227: log10_cal = 16'b0000010101000100;
            15'd21228: log10_cal = 16'b0000010101000100;
            15'd21229: log10_cal = 16'b0000010101000100;
            15'd21230: log10_cal = 16'b0000010101000100;
            15'd21231: log10_cal = 16'b0000010101000100;
            15'd21232: log10_cal = 16'b0000010101000100;
            15'd21233: log10_cal = 16'b0000010101000100;
            15'd21234: log10_cal = 16'b0000010101000100;
            15'd21235: log10_cal = 16'b0000010101000100;
            15'd21236: log10_cal = 16'b0000010101000100;
            15'd21237: log10_cal = 16'b0000010101000100;
            15'd21238: log10_cal = 16'b0000010101000100;
            15'd21239: log10_cal = 16'b0000010101000100;
            15'd21240: log10_cal = 16'b0000010101000100;
            15'd21241: log10_cal = 16'b0000010101000100;
            15'd21242: log10_cal = 16'b0000010101000100;
            15'd21243: log10_cal = 16'b0000010101000100;
            15'd21244: log10_cal = 16'b0000010101000100;
            15'd21245: log10_cal = 16'b0000010101000100;
            15'd21246: log10_cal = 16'b0000010101000100;
            15'd21247: log10_cal = 16'b0000010101000100;
            15'd21248: log10_cal = 16'b0000010101000100;
            15'd21249: log10_cal = 16'b0000010101000100;
            15'd21250: log10_cal = 16'b0000010101000100;
            15'd21251: log10_cal = 16'b0000010101000100;
            15'd21252: log10_cal = 16'b0000010101000100;
            15'd21253: log10_cal = 16'b0000010101000100;
            15'd21254: log10_cal = 16'b0000010101000100;
            15'd21255: log10_cal = 16'b0000010101000100;
            15'd21256: log10_cal = 16'b0000010101000100;
            15'd21257: log10_cal = 16'b0000010101000100;
            15'd21258: log10_cal = 16'b0000010101000100;
            15'd21259: log10_cal = 16'b0000010101000100;
            15'd21260: log10_cal = 16'b0000010101000100;
            15'd21261: log10_cal = 16'b0000010101000100;
            15'd21262: log10_cal = 16'b0000010101000100;
            15'd21263: log10_cal = 16'b0000010101000100;
            15'd21264: log10_cal = 16'b0000010101000100;
            15'd21265: log10_cal = 16'b0000010101000100;
            15'd21266: log10_cal = 16'b0000010101000101;
            15'd21267: log10_cal = 16'b0000010101000101;
            15'd21268: log10_cal = 16'b0000010101000101;
            15'd21269: log10_cal = 16'b0000010101000101;
            15'd21270: log10_cal = 16'b0000010101000101;
            15'd21271: log10_cal = 16'b0000010101000101;
            15'd21272: log10_cal = 16'b0000010101000101;
            15'd21273: log10_cal = 16'b0000010101000101;
            15'd21274: log10_cal = 16'b0000010101000101;
            15'd21275: log10_cal = 16'b0000010101000101;
            15'd21276: log10_cal = 16'b0000010101000101;
            15'd21277: log10_cal = 16'b0000010101000101;
            15'd21278: log10_cal = 16'b0000010101000101;
            15'd21279: log10_cal = 16'b0000010101000101;
            15'd21280: log10_cal = 16'b0000010101000101;
            15'd21281: log10_cal = 16'b0000010101000101;
            15'd21282: log10_cal = 16'b0000010101000101;
            15'd21283: log10_cal = 16'b0000010101000101;
            15'd21284: log10_cal = 16'b0000010101000101;
            15'd21285: log10_cal = 16'b0000010101000101;
            15'd21286: log10_cal = 16'b0000010101000101;
            15'd21287: log10_cal = 16'b0000010101000101;
            15'd21288: log10_cal = 16'b0000010101000101;
            15'd21289: log10_cal = 16'b0000010101000101;
            15'd21290: log10_cal = 16'b0000010101000101;
            15'd21291: log10_cal = 16'b0000010101000101;
            15'd21292: log10_cal = 16'b0000010101000101;
            15'd21293: log10_cal = 16'b0000010101000101;
            15'd21294: log10_cal = 16'b0000010101000101;
            15'd21295: log10_cal = 16'b0000010101000101;
            15'd21296: log10_cal = 16'b0000010101000101;
            15'd21297: log10_cal = 16'b0000010101000101;
            15'd21298: log10_cal = 16'b0000010101000101;
            15'd21299: log10_cal = 16'b0000010101000101;
            15'd21300: log10_cal = 16'b0000010101000101;
            15'd21301: log10_cal = 16'b0000010101000101;
            15'd21302: log10_cal = 16'b0000010101000101;
            15'd21303: log10_cal = 16'b0000010101000101;
            15'd21304: log10_cal = 16'b0000010101000101;
            15'd21305: log10_cal = 16'b0000010101000101;
            15'd21306: log10_cal = 16'b0000010101000101;
            15'd21307: log10_cal = 16'b0000010101000101;
            15'd21308: log10_cal = 16'b0000010101000101;
            15'd21309: log10_cal = 16'b0000010101000101;
            15'd21310: log10_cal = 16'b0000010101000101;
            15'd21311: log10_cal = 16'b0000010101000101;
            15'd21312: log10_cal = 16'b0000010101000101;
            15'd21313: log10_cal = 16'b0000010101000101;
            15'd21314: log10_cal = 16'b0000010101000110;
            15'd21315: log10_cal = 16'b0000010101000110;
            15'd21316: log10_cal = 16'b0000010101000110;
            15'd21317: log10_cal = 16'b0000010101000110;
            15'd21318: log10_cal = 16'b0000010101000110;
            15'd21319: log10_cal = 16'b0000010101000110;
            15'd21320: log10_cal = 16'b0000010101000110;
            15'd21321: log10_cal = 16'b0000010101000110;
            15'd21322: log10_cal = 16'b0000010101000110;
            15'd21323: log10_cal = 16'b0000010101000110;
            15'd21324: log10_cal = 16'b0000010101000110;
            15'd21325: log10_cal = 16'b0000010101000110;
            15'd21326: log10_cal = 16'b0000010101000110;
            15'd21327: log10_cal = 16'b0000010101000110;
            15'd21328: log10_cal = 16'b0000010101000110;
            15'd21329: log10_cal = 16'b0000010101000110;
            15'd21330: log10_cal = 16'b0000010101000110;
            15'd21331: log10_cal = 16'b0000010101000110;
            15'd21332: log10_cal = 16'b0000010101000110;
            15'd21333: log10_cal = 16'b0000010101000110;
            15'd21334: log10_cal = 16'b0000010101000110;
            15'd21335: log10_cal = 16'b0000010101000110;
            15'd21336: log10_cal = 16'b0000010101000110;
            15'd21337: log10_cal = 16'b0000010101000110;
            15'd21338: log10_cal = 16'b0000010101000110;
            15'd21339: log10_cal = 16'b0000010101000110;
            15'd21340: log10_cal = 16'b0000010101000110;
            15'd21341: log10_cal = 16'b0000010101000110;
            15'd21342: log10_cal = 16'b0000010101000110;
            15'd21343: log10_cal = 16'b0000010101000110;
            15'd21344: log10_cal = 16'b0000010101000110;
            15'd21345: log10_cal = 16'b0000010101000110;
            15'd21346: log10_cal = 16'b0000010101000110;
            15'd21347: log10_cal = 16'b0000010101000110;
            15'd21348: log10_cal = 16'b0000010101000110;
            15'd21349: log10_cal = 16'b0000010101000110;
            15'd21350: log10_cal = 16'b0000010101000110;
            15'd21351: log10_cal = 16'b0000010101000110;
            15'd21352: log10_cal = 16'b0000010101000110;
            15'd21353: log10_cal = 16'b0000010101000110;
            15'd21354: log10_cal = 16'b0000010101000110;
            15'd21355: log10_cal = 16'b0000010101000110;
            15'd21356: log10_cal = 16'b0000010101000110;
            15'd21357: log10_cal = 16'b0000010101000110;
            15'd21358: log10_cal = 16'b0000010101000110;
            15'd21359: log10_cal = 16'b0000010101000110;
            15'd21360: log10_cal = 16'b0000010101000110;
            15'd21361: log10_cal = 16'b0000010101000110;
            15'd21362: log10_cal = 16'b0000010101000111;
            15'd21363: log10_cal = 16'b0000010101000111;
            15'd21364: log10_cal = 16'b0000010101000111;
            15'd21365: log10_cal = 16'b0000010101000111;
            15'd21366: log10_cal = 16'b0000010101000111;
            15'd21367: log10_cal = 16'b0000010101000111;
            15'd21368: log10_cal = 16'b0000010101000111;
            15'd21369: log10_cal = 16'b0000010101000111;
            15'd21370: log10_cal = 16'b0000010101000111;
            15'd21371: log10_cal = 16'b0000010101000111;
            15'd21372: log10_cal = 16'b0000010101000111;
            15'd21373: log10_cal = 16'b0000010101000111;
            15'd21374: log10_cal = 16'b0000010101000111;
            15'd21375: log10_cal = 16'b0000010101000111;
            15'd21376: log10_cal = 16'b0000010101000111;
            15'd21377: log10_cal = 16'b0000010101000111;
            15'd21378: log10_cal = 16'b0000010101000111;
            15'd21379: log10_cal = 16'b0000010101000111;
            15'd21380: log10_cal = 16'b0000010101000111;
            15'd21381: log10_cal = 16'b0000010101000111;
            15'd21382: log10_cal = 16'b0000010101000111;
            15'd21383: log10_cal = 16'b0000010101000111;
            15'd21384: log10_cal = 16'b0000010101000111;
            15'd21385: log10_cal = 16'b0000010101000111;
            15'd21386: log10_cal = 16'b0000010101000111;
            15'd21387: log10_cal = 16'b0000010101000111;
            15'd21388: log10_cal = 16'b0000010101000111;
            15'd21389: log10_cal = 16'b0000010101000111;
            15'd21390: log10_cal = 16'b0000010101000111;
            15'd21391: log10_cal = 16'b0000010101000111;
            15'd21392: log10_cal = 16'b0000010101000111;
            15'd21393: log10_cal = 16'b0000010101000111;
            15'd21394: log10_cal = 16'b0000010101000111;
            15'd21395: log10_cal = 16'b0000010101000111;
            15'd21396: log10_cal = 16'b0000010101000111;
            15'd21397: log10_cal = 16'b0000010101000111;
            15'd21398: log10_cal = 16'b0000010101000111;
            15'd21399: log10_cal = 16'b0000010101000111;
            15'd21400: log10_cal = 16'b0000010101000111;
            15'd21401: log10_cal = 16'b0000010101000111;
            15'd21402: log10_cal = 16'b0000010101000111;
            15'd21403: log10_cal = 16'b0000010101000111;
            15'd21404: log10_cal = 16'b0000010101000111;
            15'd21405: log10_cal = 16'b0000010101000111;
            15'd21406: log10_cal = 16'b0000010101000111;
            15'd21407: log10_cal = 16'b0000010101000111;
            15'd21408: log10_cal = 16'b0000010101000111;
            15'd21409: log10_cal = 16'b0000010101000111;
            15'd21410: log10_cal = 16'b0000010101001000;
            15'd21411: log10_cal = 16'b0000010101001000;
            15'd21412: log10_cal = 16'b0000010101001000;
            15'd21413: log10_cal = 16'b0000010101001000;
            15'd21414: log10_cal = 16'b0000010101001000;
            15'd21415: log10_cal = 16'b0000010101001000;
            15'd21416: log10_cal = 16'b0000010101001000;
            15'd21417: log10_cal = 16'b0000010101001000;
            15'd21418: log10_cal = 16'b0000010101001000;
            15'd21419: log10_cal = 16'b0000010101001000;
            15'd21420: log10_cal = 16'b0000010101001000;
            15'd21421: log10_cal = 16'b0000010101001000;
            15'd21422: log10_cal = 16'b0000010101001000;
            15'd21423: log10_cal = 16'b0000010101001000;
            15'd21424: log10_cal = 16'b0000010101001000;
            15'd21425: log10_cal = 16'b0000010101001000;
            15'd21426: log10_cal = 16'b0000010101001000;
            15'd21427: log10_cal = 16'b0000010101001000;
            15'd21428: log10_cal = 16'b0000010101001000;
            15'd21429: log10_cal = 16'b0000010101001000;
            15'd21430: log10_cal = 16'b0000010101001000;
            15'd21431: log10_cal = 16'b0000010101001000;
            15'd21432: log10_cal = 16'b0000010101001000;
            15'd21433: log10_cal = 16'b0000010101001000;
            15'd21434: log10_cal = 16'b0000010101001000;
            15'd21435: log10_cal = 16'b0000010101001000;
            15'd21436: log10_cal = 16'b0000010101001000;
            15'd21437: log10_cal = 16'b0000010101001000;
            15'd21438: log10_cal = 16'b0000010101001000;
            15'd21439: log10_cal = 16'b0000010101001000;
            15'd21440: log10_cal = 16'b0000010101001000;
            15'd21441: log10_cal = 16'b0000010101001000;
            15'd21442: log10_cal = 16'b0000010101001000;
            15'd21443: log10_cal = 16'b0000010101001000;
            15'd21444: log10_cal = 16'b0000010101001000;
            15'd21445: log10_cal = 16'b0000010101001000;
            15'd21446: log10_cal = 16'b0000010101001000;
            15'd21447: log10_cal = 16'b0000010101001000;
            15'd21448: log10_cal = 16'b0000010101001000;
            15'd21449: log10_cal = 16'b0000010101001000;
            15'd21450: log10_cal = 16'b0000010101001000;
            15'd21451: log10_cal = 16'b0000010101001000;
            15'd21452: log10_cal = 16'b0000010101001000;
            15'd21453: log10_cal = 16'b0000010101001000;
            15'd21454: log10_cal = 16'b0000010101001000;
            15'd21455: log10_cal = 16'b0000010101001000;
            15'd21456: log10_cal = 16'b0000010101001000;
            15'd21457: log10_cal = 16'b0000010101001000;
            15'd21458: log10_cal = 16'b0000010101001001;
            15'd21459: log10_cal = 16'b0000010101001001;
            15'd21460: log10_cal = 16'b0000010101001001;
            15'd21461: log10_cal = 16'b0000010101001001;
            15'd21462: log10_cal = 16'b0000010101001001;
            15'd21463: log10_cal = 16'b0000010101001001;
            15'd21464: log10_cal = 16'b0000010101001001;
            15'd21465: log10_cal = 16'b0000010101001001;
            15'd21466: log10_cal = 16'b0000010101001001;
            15'd21467: log10_cal = 16'b0000010101001001;
            15'd21468: log10_cal = 16'b0000010101001001;
            15'd21469: log10_cal = 16'b0000010101001001;
            15'd21470: log10_cal = 16'b0000010101001001;
            15'd21471: log10_cal = 16'b0000010101001001;
            15'd21472: log10_cal = 16'b0000010101001001;
            15'd21473: log10_cal = 16'b0000010101001001;
            15'd21474: log10_cal = 16'b0000010101001001;
            15'd21475: log10_cal = 16'b0000010101001001;
            15'd21476: log10_cal = 16'b0000010101001001;
            15'd21477: log10_cal = 16'b0000010101001001;
            15'd21478: log10_cal = 16'b0000010101001001;
            15'd21479: log10_cal = 16'b0000010101001001;
            15'd21480: log10_cal = 16'b0000010101001001;
            15'd21481: log10_cal = 16'b0000010101001001;
            15'd21482: log10_cal = 16'b0000010101001001;
            15'd21483: log10_cal = 16'b0000010101001001;
            15'd21484: log10_cal = 16'b0000010101001001;
            15'd21485: log10_cal = 16'b0000010101001001;
            15'd21486: log10_cal = 16'b0000010101001001;
            15'd21487: log10_cal = 16'b0000010101001001;
            15'd21488: log10_cal = 16'b0000010101001001;
            15'd21489: log10_cal = 16'b0000010101001001;
            15'd21490: log10_cal = 16'b0000010101001001;
            15'd21491: log10_cal = 16'b0000010101001001;
            15'd21492: log10_cal = 16'b0000010101001001;
            15'd21493: log10_cal = 16'b0000010101001001;
            15'd21494: log10_cal = 16'b0000010101001001;
            15'd21495: log10_cal = 16'b0000010101001001;
            15'd21496: log10_cal = 16'b0000010101001001;
            15'd21497: log10_cal = 16'b0000010101001001;
            15'd21498: log10_cal = 16'b0000010101001001;
            15'd21499: log10_cal = 16'b0000010101001001;
            15'd21500: log10_cal = 16'b0000010101001001;
            15'd21501: log10_cal = 16'b0000010101001001;
            15'd21502: log10_cal = 16'b0000010101001001;
            15'd21503: log10_cal = 16'b0000010101001001;
            15'd21504: log10_cal = 16'b0000010101001001;
            15'd21505: log10_cal = 16'b0000010101001001;
            15'd21506: log10_cal = 16'b0000010101001001;
            15'd21507: log10_cal = 16'b0000010101001010;
            15'd21508: log10_cal = 16'b0000010101001010;
            15'd21509: log10_cal = 16'b0000010101001010;
            15'd21510: log10_cal = 16'b0000010101001010;
            15'd21511: log10_cal = 16'b0000010101001010;
            15'd21512: log10_cal = 16'b0000010101001010;
            15'd21513: log10_cal = 16'b0000010101001010;
            15'd21514: log10_cal = 16'b0000010101001010;
            15'd21515: log10_cal = 16'b0000010101001010;
            15'd21516: log10_cal = 16'b0000010101001010;
            15'd21517: log10_cal = 16'b0000010101001010;
            15'd21518: log10_cal = 16'b0000010101001010;
            15'd21519: log10_cal = 16'b0000010101001010;
            15'd21520: log10_cal = 16'b0000010101001010;
            15'd21521: log10_cal = 16'b0000010101001010;
            15'd21522: log10_cal = 16'b0000010101001010;
            15'd21523: log10_cal = 16'b0000010101001010;
            15'd21524: log10_cal = 16'b0000010101001010;
            15'd21525: log10_cal = 16'b0000010101001010;
            15'd21526: log10_cal = 16'b0000010101001010;
            15'd21527: log10_cal = 16'b0000010101001010;
            15'd21528: log10_cal = 16'b0000010101001010;
            15'd21529: log10_cal = 16'b0000010101001010;
            15'd21530: log10_cal = 16'b0000010101001010;
            15'd21531: log10_cal = 16'b0000010101001010;
            15'd21532: log10_cal = 16'b0000010101001010;
            15'd21533: log10_cal = 16'b0000010101001010;
            15'd21534: log10_cal = 16'b0000010101001010;
            15'd21535: log10_cal = 16'b0000010101001010;
            15'd21536: log10_cal = 16'b0000010101001010;
            15'd21537: log10_cal = 16'b0000010101001010;
            15'd21538: log10_cal = 16'b0000010101001010;
            15'd21539: log10_cal = 16'b0000010101001010;
            15'd21540: log10_cal = 16'b0000010101001010;
            15'd21541: log10_cal = 16'b0000010101001010;
            15'd21542: log10_cal = 16'b0000010101001010;
            15'd21543: log10_cal = 16'b0000010101001010;
            15'd21544: log10_cal = 16'b0000010101001010;
            15'd21545: log10_cal = 16'b0000010101001010;
            15'd21546: log10_cal = 16'b0000010101001010;
            15'd21547: log10_cal = 16'b0000010101001010;
            15'd21548: log10_cal = 16'b0000010101001010;
            15'd21549: log10_cal = 16'b0000010101001010;
            15'd21550: log10_cal = 16'b0000010101001010;
            15'd21551: log10_cal = 16'b0000010101001010;
            15'd21552: log10_cal = 16'b0000010101001010;
            15'd21553: log10_cal = 16'b0000010101001010;
            15'd21554: log10_cal = 16'b0000010101001010;
            15'd21555: log10_cal = 16'b0000010101001011;
            15'd21556: log10_cal = 16'b0000010101001011;
            15'd21557: log10_cal = 16'b0000010101001011;
            15'd21558: log10_cal = 16'b0000010101001011;
            15'd21559: log10_cal = 16'b0000010101001011;
            15'd21560: log10_cal = 16'b0000010101001011;
            15'd21561: log10_cal = 16'b0000010101001011;
            15'd21562: log10_cal = 16'b0000010101001011;
            15'd21563: log10_cal = 16'b0000010101001011;
            15'd21564: log10_cal = 16'b0000010101001011;
            15'd21565: log10_cal = 16'b0000010101001011;
            15'd21566: log10_cal = 16'b0000010101001011;
            15'd21567: log10_cal = 16'b0000010101001011;
            15'd21568: log10_cal = 16'b0000010101001011;
            15'd21569: log10_cal = 16'b0000010101001011;
            15'd21570: log10_cal = 16'b0000010101001011;
            15'd21571: log10_cal = 16'b0000010101001011;
            15'd21572: log10_cal = 16'b0000010101001011;
            15'd21573: log10_cal = 16'b0000010101001011;
            15'd21574: log10_cal = 16'b0000010101001011;
            15'd21575: log10_cal = 16'b0000010101001011;
            15'd21576: log10_cal = 16'b0000010101001011;
            15'd21577: log10_cal = 16'b0000010101001011;
            15'd21578: log10_cal = 16'b0000010101001011;
            15'd21579: log10_cal = 16'b0000010101001011;
            15'd21580: log10_cal = 16'b0000010101001011;
            15'd21581: log10_cal = 16'b0000010101001011;
            15'd21582: log10_cal = 16'b0000010101001011;
            15'd21583: log10_cal = 16'b0000010101001011;
            15'd21584: log10_cal = 16'b0000010101001011;
            15'd21585: log10_cal = 16'b0000010101001011;
            15'd21586: log10_cal = 16'b0000010101001011;
            15'd21587: log10_cal = 16'b0000010101001011;
            15'd21588: log10_cal = 16'b0000010101001011;
            15'd21589: log10_cal = 16'b0000010101001011;
            15'd21590: log10_cal = 16'b0000010101001011;
            15'd21591: log10_cal = 16'b0000010101001011;
            15'd21592: log10_cal = 16'b0000010101001011;
            15'd21593: log10_cal = 16'b0000010101001011;
            15'd21594: log10_cal = 16'b0000010101001011;
            15'd21595: log10_cal = 16'b0000010101001011;
            15'd21596: log10_cal = 16'b0000010101001011;
            15'd21597: log10_cal = 16'b0000010101001011;
            15'd21598: log10_cal = 16'b0000010101001011;
            15'd21599: log10_cal = 16'b0000010101001011;
            15'd21600: log10_cal = 16'b0000010101001011;
            15'd21601: log10_cal = 16'b0000010101001011;
            15'd21602: log10_cal = 16'b0000010101001011;
            15'd21603: log10_cal = 16'b0000010101001011;
            15'd21604: log10_cal = 16'b0000010101001100;
            15'd21605: log10_cal = 16'b0000010101001100;
            15'd21606: log10_cal = 16'b0000010101001100;
            15'd21607: log10_cal = 16'b0000010101001100;
            15'd21608: log10_cal = 16'b0000010101001100;
            15'd21609: log10_cal = 16'b0000010101001100;
            15'd21610: log10_cal = 16'b0000010101001100;
            15'd21611: log10_cal = 16'b0000010101001100;
            15'd21612: log10_cal = 16'b0000010101001100;
            15'd21613: log10_cal = 16'b0000010101001100;
            15'd21614: log10_cal = 16'b0000010101001100;
            15'd21615: log10_cal = 16'b0000010101001100;
            15'd21616: log10_cal = 16'b0000010101001100;
            15'd21617: log10_cal = 16'b0000010101001100;
            15'd21618: log10_cal = 16'b0000010101001100;
            15'd21619: log10_cal = 16'b0000010101001100;
            15'd21620: log10_cal = 16'b0000010101001100;
            15'd21621: log10_cal = 16'b0000010101001100;
            15'd21622: log10_cal = 16'b0000010101001100;
            15'd21623: log10_cal = 16'b0000010101001100;
            15'd21624: log10_cal = 16'b0000010101001100;
            15'd21625: log10_cal = 16'b0000010101001100;
            15'd21626: log10_cal = 16'b0000010101001100;
            15'd21627: log10_cal = 16'b0000010101001100;
            15'd21628: log10_cal = 16'b0000010101001100;
            15'd21629: log10_cal = 16'b0000010101001100;
            15'd21630: log10_cal = 16'b0000010101001100;
            15'd21631: log10_cal = 16'b0000010101001100;
            15'd21632: log10_cal = 16'b0000010101001100;
            15'd21633: log10_cal = 16'b0000010101001100;
            15'd21634: log10_cal = 16'b0000010101001100;
            15'd21635: log10_cal = 16'b0000010101001100;
            15'd21636: log10_cal = 16'b0000010101001100;
            15'd21637: log10_cal = 16'b0000010101001100;
            15'd21638: log10_cal = 16'b0000010101001100;
            15'd21639: log10_cal = 16'b0000010101001100;
            15'd21640: log10_cal = 16'b0000010101001100;
            15'd21641: log10_cal = 16'b0000010101001100;
            15'd21642: log10_cal = 16'b0000010101001100;
            15'd21643: log10_cal = 16'b0000010101001100;
            15'd21644: log10_cal = 16'b0000010101001100;
            15'd21645: log10_cal = 16'b0000010101001100;
            15'd21646: log10_cal = 16'b0000010101001100;
            15'd21647: log10_cal = 16'b0000010101001100;
            15'd21648: log10_cal = 16'b0000010101001100;
            15'd21649: log10_cal = 16'b0000010101001100;
            15'd21650: log10_cal = 16'b0000010101001100;
            15'd21651: log10_cal = 16'b0000010101001100;
            15'd21652: log10_cal = 16'b0000010101001101;
            15'd21653: log10_cal = 16'b0000010101001101;
            15'd21654: log10_cal = 16'b0000010101001101;
            15'd21655: log10_cal = 16'b0000010101001101;
            15'd21656: log10_cal = 16'b0000010101001101;
            15'd21657: log10_cal = 16'b0000010101001101;
            15'd21658: log10_cal = 16'b0000010101001101;
            15'd21659: log10_cal = 16'b0000010101001101;
            15'd21660: log10_cal = 16'b0000010101001101;
            15'd21661: log10_cal = 16'b0000010101001101;
            15'd21662: log10_cal = 16'b0000010101001101;
            15'd21663: log10_cal = 16'b0000010101001101;
            15'd21664: log10_cal = 16'b0000010101001101;
            15'd21665: log10_cal = 16'b0000010101001101;
            15'd21666: log10_cal = 16'b0000010101001101;
            15'd21667: log10_cal = 16'b0000010101001101;
            15'd21668: log10_cal = 16'b0000010101001101;
            15'd21669: log10_cal = 16'b0000010101001101;
            15'd21670: log10_cal = 16'b0000010101001101;
            15'd21671: log10_cal = 16'b0000010101001101;
            15'd21672: log10_cal = 16'b0000010101001101;
            15'd21673: log10_cal = 16'b0000010101001101;
            15'd21674: log10_cal = 16'b0000010101001101;
            15'd21675: log10_cal = 16'b0000010101001101;
            15'd21676: log10_cal = 16'b0000010101001101;
            15'd21677: log10_cal = 16'b0000010101001101;
            15'd21678: log10_cal = 16'b0000010101001101;
            15'd21679: log10_cal = 16'b0000010101001101;
            15'd21680: log10_cal = 16'b0000010101001101;
            15'd21681: log10_cal = 16'b0000010101001101;
            15'd21682: log10_cal = 16'b0000010101001101;
            15'd21683: log10_cal = 16'b0000010101001101;
            15'd21684: log10_cal = 16'b0000010101001101;
            15'd21685: log10_cal = 16'b0000010101001101;
            15'd21686: log10_cal = 16'b0000010101001101;
            15'd21687: log10_cal = 16'b0000010101001101;
            15'd21688: log10_cal = 16'b0000010101001101;
            15'd21689: log10_cal = 16'b0000010101001101;
            15'd21690: log10_cal = 16'b0000010101001101;
            15'd21691: log10_cal = 16'b0000010101001101;
            15'd21692: log10_cal = 16'b0000010101001101;
            15'd21693: log10_cal = 16'b0000010101001101;
            15'd21694: log10_cal = 16'b0000010101001101;
            15'd21695: log10_cal = 16'b0000010101001101;
            15'd21696: log10_cal = 16'b0000010101001101;
            15'd21697: log10_cal = 16'b0000010101001101;
            15'd21698: log10_cal = 16'b0000010101001101;
            15'd21699: log10_cal = 16'b0000010101001101;
            15'd21700: log10_cal = 16'b0000010101001101;
            15'd21701: log10_cal = 16'b0000010101001110;
            15'd21702: log10_cal = 16'b0000010101001110;
            15'd21703: log10_cal = 16'b0000010101001110;
            15'd21704: log10_cal = 16'b0000010101001110;
            15'd21705: log10_cal = 16'b0000010101001110;
            15'd21706: log10_cal = 16'b0000010101001110;
            15'd21707: log10_cal = 16'b0000010101001110;
            15'd21708: log10_cal = 16'b0000010101001110;
            15'd21709: log10_cal = 16'b0000010101001110;
            15'd21710: log10_cal = 16'b0000010101001110;
            15'd21711: log10_cal = 16'b0000010101001110;
            15'd21712: log10_cal = 16'b0000010101001110;
            15'd21713: log10_cal = 16'b0000010101001110;
            15'd21714: log10_cal = 16'b0000010101001110;
            15'd21715: log10_cal = 16'b0000010101001110;
            15'd21716: log10_cal = 16'b0000010101001110;
            15'd21717: log10_cal = 16'b0000010101001110;
            15'd21718: log10_cal = 16'b0000010101001110;
            15'd21719: log10_cal = 16'b0000010101001110;
            15'd21720: log10_cal = 16'b0000010101001110;
            15'd21721: log10_cal = 16'b0000010101001110;
            15'd21722: log10_cal = 16'b0000010101001110;
            15'd21723: log10_cal = 16'b0000010101001110;
            15'd21724: log10_cal = 16'b0000010101001110;
            15'd21725: log10_cal = 16'b0000010101001110;
            15'd21726: log10_cal = 16'b0000010101001110;
            15'd21727: log10_cal = 16'b0000010101001110;
            15'd21728: log10_cal = 16'b0000010101001110;
            15'd21729: log10_cal = 16'b0000010101001110;
            15'd21730: log10_cal = 16'b0000010101001110;
            15'd21731: log10_cal = 16'b0000010101001110;
            15'd21732: log10_cal = 16'b0000010101001110;
            15'd21733: log10_cal = 16'b0000010101001110;
            15'd21734: log10_cal = 16'b0000010101001110;
            15'd21735: log10_cal = 16'b0000010101001110;
            15'd21736: log10_cal = 16'b0000010101001110;
            15'd21737: log10_cal = 16'b0000010101001110;
            15'd21738: log10_cal = 16'b0000010101001110;
            15'd21739: log10_cal = 16'b0000010101001110;
            15'd21740: log10_cal = 16'b0000010101001110;
            15'd21741: log10_cal = 16'b0000010101001110;
            15'd21742: log10_cal = 16'b0000010101001110;
            15'd21743: log10_cal = 16'b0000010101001110;
            15'd21744: log10_cal = 16'b0000010101001110;
            15'd21745: log10_cal = 16'b0000010101001110;
            15'd21746: log10_cal = 16'b0000010101001110;
            15'd21747: log10_cal = 16'b0000010101001110;
            15'd21748: log10_cal = 16'b0000010101001110;
            15'd21749: log10_cal = 16'b0000010101001110;
            15'd21750: log10_cal = 16'b0000010101001111;
            15'd21751: log10_cal = 16'b0000010101001111;
            15'd21752: log10_cal = 16'b0000010101001111;
            15'd21753: log10_cal = 16'b0000010101001111;
            15'd21754: log10_cal = 16'b0000010101001111;
            15'd21755: log10_cal = 16'b0000010101001111;
            15'd21756: log10_cal = 16'b0000010101001111;
            15'd21757: log10_cal = 16'b0000010101001111;
            15'd21758: log10_cal = 16'b0000010101001111;
            15'd21759: log10_cal = 16'b0000010101001111;
            15'd21760: log10_cal = 16'b0000010101001111;
            15'd21761: log10_cal = 16'b0000010101001111;
            15'd21762: log10_cal = 16'b0000010101001111;
            15'd21763: log10_cal = 16'b0000010101001111;
            15'd21764: log10_cal = 16'b0000010101001111;
            15'd21765: log10_cal = 16'b0000010101001111;
            15'd21766: log10_cal = 16'b0000010101001111;
            15'd21767: log10_cal = 16'b0000010101001111;
            15'd21768: log10_cal = 16'b0000010101001111;
            15'd21769: log10_cal = 16'b0000010101001111;
            15'd21770: log10_cal = 16'b0000010101001111;
            15'd21771: log10_cal = 16'b0000010101001111;
            15'd21772: log10_cal = 16'b0000010101001111;
            15'd21773: log10_cal = 16'b0000010101001111;
            15'd21774: log10_cal = 16'b0000010101001111;
            15'd21775: log10_cal = 16'b0000010101001111;
            15'd21776: log10_cal = 16'b0000010101001111;
            15'd21777: log10_cal = 16'b0000010101001111;
            15'd21778: log10_cal = 16'b0000010101001111;
            15'd21779: log10_cal = 16'b0000010101001111;
            15'd21780: log10_cal = 16'b0000010101001111;
            15'd21781: log10_cal = 16'b0000010101001111;
            15'd21782: log10_cal = 16'b0000010101001111;
            15'd21783: log10_cal = 16'b0000010101001111;
            15'd21784: log10_cal = 16'b0000010101001111;
            15'd21785: log10_cal = 16'b0000010101001111;
            15'd21786: log10_cal = 16'b0000010101001111;
            15'd21787: log10_cal = 16'b0000010101001111;
            15'd21788: log10_cal = 16'b0000010101001111;
            15'd21789: log10_cal = 16'b0000010101001111;
            15'd21790: log10_cal = 16'b0000010101001111;
            15'd21791: log10_cal = 16'b0000010101001111;
            15'd21792: log10_cal = 16'b0000010101001111;
            15'd21793: log10_cal = 16'b0000010101001111;
            15'd21794: log10_cal = 16'b0000010101001111;
            15'd21795: log10_cal = 16'b0000010101001111;
            15'd21796: log10_cal = 16'b0000010101001111;
            15'd21797: log10_cal = 16'b0000010101001111;
            15'd21798: log10_cal = 16'b0000010101001111;
            15'd21799: log10_cal = 16'b0000010101010000;
            15'd21800: log10_cal = 16'b0000010101010000;
            15'd21801: log10_cal = 16'b0000010101010000;
            15'd21802: log10_cal = 16'b0000010101010000;
            15'd21803: log10_cal = 16'b0000010101010000;
            15'd21804: log10_cal = 16'b0000010101010000;
            15'd21805: log10_cal = 16'b0000010101010000;
            15'd21806: log10_cal = 16'b0000010101010000;
            15'd21807: log10_cal = 16'b0000010101010000;
            15'd21808: log10_cal = 16'b0000010101010000;
            15'd21809: log10_cal = 16'b0000010101010000;
            15'd21810: log10_cal = 16'b0000010101010000;
            15'd21811: log10_cal = 16'b0000010101010000;
            15'd21812: log10_cal = 16'b0000010101010000;
            15'd21813: log10_cal = 16'b0000010101010000;
            15'd21814: log10_cal = 16'b0000010101010000;
            15'd21815: log10_cal = 16'b0000010101010000;
            15'd21816: log10_cal = 16'b0000010101010000;
            15'd21817: log10_cal = 16'b0000010101010000;
            15'd21818: log10_cal = 16'b0000010101010000;
            15'd21819: log10_cal = 16'b0000010101010000;
            15'd21820: log10_cal = 16'b0000010101010000;
            15'd21821: log10_cal = 16'b0000010101010000;
            15'd21822: log10_cal = 16'b0000010101010000;
            15'd21823: log10_cal = 16'b0000010101010000;
            15'd21824: log10_cal = 16'b0000010101010000;
            15'd21825: log10_cal = 16'b0000010101010000;
            15'd21826: log10_cal = 16'b0000010101010000;
            15'd21827: log10_cal = 16'b0000010101010000;
            15'd21828: log10_cal = 16'b0000010101010000;
            15'd21829: log10_cal = 16'b0000010101010000;
            15'd21830: log10_cal = 16'b0000010101010000;
            15'd21831: log10_cal = 16'b0000010101010000;
            15'd21832: log10_cal = 16'b0000010101010000;
            15'd21833: log10_cal = 16'b0000010101010000;
            15'd21834: log10_cal = 16'b0000010101010000;
            15'd21835: log10_cal = 16'b0000010101010000;
            15'd21836: log10_cal = 16'b0000010101010000;
            15'd21837: log10_cal = 16'b0000010101010000;
            15'd21838: log10_cal = 16'b0000010101010000;
            15'd21839: log10_cal = 16'b0000010101010000;
            15'd21840: log10_cal = 16'b0000010101010000;
            15'd21841: log10_cal = 16'b0000010101010000;
            15'd21842: log10_cal = 16'b0000010101010000;
            15'd21843: log10_cal = 16'b0000010101010000;
            15'd21844: log10_cal = 16'b0000010101010000;
            15'd21845: log10_cal = 16'b0000010101010000;
            15'd21846: log10_cal = 16'b0000010101010000;
            15'd21847: log10_cal = 16'b0000010101010000;
            15'd21848: log10_cal = 16'b0000010101010001;
            15'd21849: log10_cal = 16'b0000010101010001;
            15'd21850: log10_cal = 16'b0000010101010001;
            15'd21851: log10_cal = 16'b0000010101010001;
            15'd21852: log10_cal = 16'b0000010101010001;
            15'd21853: log10_cal = 16'b0000010101010001;
            15'd21854: log10_cal = 16'b0000010101010001;
            15'd21855: log10_cal = 16'b0000010101010001;
            15'd21856: log10_cal = 16'b0000010101010001;
            15'd21857: log10_cal = 16'b0000010101010001;
            15'd21858: log10_cal = 16'b0000010101010001;
            15'd21859: log10_cal = 16'b0000010101010001;
            15'd21860: log10_cal = 16'b0000010101010001;
            15'd21861: log10_cal = 16'b0000010101010001;
            15'd21862: log10_cal = 16'b0000010101010001;
            15'd21863: log10_cal = 16'b0000010101010001;
            15'd21864: log10_cal = 16'b0000010101010001;
            15'd21865: log10_cal = 16'b0000010101010001;
            15'd21866: log10_cal = 16'b0000010101010001;
            15'd21867: log10_cal = 16'b0000010101010001;
            15'd21868: log10_cal = 16'b0000010101010001;
            15'd21869: log10_cal = 16'b0000010101010001;
            15'd21870: log10_cal = 16'b0000010101010001;
            15'd21871: log10_cal = 16'b0000010101010001;
            15'd21872: log10_cal = 16'b0000010101010001;
            15'd21873: log10_cal = 16'b0000010101010001;
            15'd21874: log10_cal = 16'b0000010101010001;
            15'd21875: log10_cal = 16'b0000010101010001;
            15'd21876: log10_cal = 16'b0000010101010001;
            15'd21877: log10_cal = 16'b0000010101010001;
            15'd21878: log10_cal = 16'b0000010101010001;
            15'd21879: log10_cal = 16'b0000010101010001;
            15'd21880: log10_cal = 16'b0000010101010001;
            15'd21881: log10_cal = 16'b0000010101010001;
            15'd21882: log10_cal = 16'b0000010101010001;
            15'd21883: log10_cal = 16'b0000010101010001;
            15'd21884: log10_cal = 16'b0000010101010001;
            15'd21885: log10_cal = 16'b0000010101010001;
            15'd21886: log10_cal = 16'b0000010101010001;
            15'd21887: log10_cal = 16'b0000010101010001;
            15'd21888: log10_cal = 16'b0000010101010001;
            15'd21889: log10_cal = 16'b0000010101010001;
            15'd21890: log10_cal = 16'b0000010101010001;
            15'd21891: log10_cal = 16'b0000010101010001;
            15'd21892: log10_cal = 16'b0000010101010001;
            15'd21893: log10_cal = 16'b0000010101010001;
            15'd21894: log10_cal = 16'b0000010101010001;
            15'd21895: log10_cal = 16'b0000010101010001;
            15'd21896: log10_cal = 16'b0000010101010001;
            15'd21897: log10_cal = 16'b0000010101010010;
            15'd21898: log10_cal = 16'b0000010101010010;
            15'd21899: log10_cal = 16'b0000010101010010;
            15'd21900: log10_cal = 16'b0000010101010010;
            15'd21901: log10_cal = 16'b0000010101010010;
            15'd21902: log10_cal = 16'b0000010101010010;
            15'd21903: log10_cal = 16'b0000010101010010;
            15'd21904: log10_cal = 16'b0000010101010010;
            15'd21905: log10_cal = 16'b0000010101010010;
            15'd21906: log10_cal = 16'b0000010101010010;
            15'd21907: log10_cal = 16'b0000010101010010;
            15'd21908: log10_cal = 16'b0000010101010010;
            15'd21909: log10_cal = 16'b0000010101010010;
            15'd21910: log10_cal = 16'b0000010101010010;
            15'd21911: log10_cal = 16'b0000010101010010;
            15'd21912: log10_cal = 16'b0000010101010010;
            15'd21913: log10_cal = 16'b0000010101010010;
            15'd21914: log10_cal = 16'b0000010101010010;
            15'd21915: log10_cal = 16'b0000010101010010;
            15'd21916: log10_cal = 16'b0000010101010010;
            15'd21917: log10_cal = 16'b0000010101010010;
            15'd21918: log10_cal = 16'b0000010101010010;
            15'd21919: log10_cal = 16'b0000010101010010;
            15'd21920: log10_cal = 16'b0000010101010010;
            15'd21921: log10_cal = 16'b0000010101010010;
            15'd21922: log10_cal = 16'b0000010101010010;
            15'd21923: log10_cal = 16'b0000010101010010;
            15'd21924: log10_cal = 16'b0000010101010010;
            15'd21925: log10_cal = 16'b0000010101010010;
            15'd21926: log10_cal = 16'b0000010101010010;
            15'd21927: log10_cal = 16'b0000010101010010;
            15'd21928: log10_cal = 16'b0000010101010010;
            15'd21929: log10_cal = 16'b0000010101010010;
            15'd21930: log10_cal = 16'b0000010101010010;
            15'd21931: log10_cal = 16'b0000010101010010;
            15'd21932: log10_cal = 16'b0000010101010010;
            15'd21933: log10_cal = 16'b0000010101010010;
            15'd21934: log10_cal = 16'b0000010101010010;
            15'd21935: log10_cal = 16'b0000010101010010;
            15'd21936: log10_cal = 16'b0000010101010010;
            15'd21937: log10_cal = 16'b0000010101010010;
            15'd21938: log10_cal = 16'b0000010101010010;
            15'd21939: log10_cal = 16'b0000010101010010;
            15'd21940: log10_cal = 16'b0000010101010010;
            15'd21941: log10_cal = 16'b0000010101010010;
            15'd21942: log10_cal = 16'b0000010101010010;
            15'd21943: log10_cal = 16'b0000010101010010;
            15'd21944: log10_cal = 16'b0000010101010010;
            15'd21945: log10_cal = 16'b0000010101010010;
            15'd21946: log10_cal = 16'b0000010101010011;
            15'd21947: log10_cal = 16'b0000010101010011;
            15'd21948: log10_cal = 16'b0000010101010011;
            15'd21949: log10_cal = 16'b0000010101010011;
            15'd21950: log10_cal = 16'b0000010101010011;
            15'd21951: log10_cal = 16'b0000010101010011;
            15'd21952: log10_cal = 16'b0000010101010011;
            15'd21953: log10_cal = 16'b0000010101010011;
            15'd21954: log10_cal = 16'b0000010101010011;
            15'd21955: log10_cal = 16'b0000010101010011;
            15'd21956: log10_cal = 16'b0000010101010011;
            15'd21957: log10_cal = 16'b0000010101010011;
            15'd21958: log10_cal = 16'b0000010101010011;
            15'd21959: log10_cal = 16'b0000010101010011;
            15'd21960: log10_cal = 16'b0000010101010011;
            15'd21961: log10_cal = 16'b0000010101010011;
            15'd21962: log10_cal = 16'b0000010101010011;
            15'd21963: log10_cal = 16'b0000010101010011;
            15'd21964: log10_cal = 16'b0000010101010011;
            15'd21965: log10_cal = 16'b0000010101010011;
            15'd21966: log10_cal = 16'b0000010101010011;
            15'd21967: log10_cal = 16'b0000010101010011;
            15'd21968: log10_cal = 16'b0000010101010011;
            15'd21969: log10_cal = 16'b0000010101010011;
            15'd21970: log10_cal = 16'b0000010101010011;
            15'd21971: log10_cal = 16'b0000010101010011;
            15'd21972: log10_cal = 16'b0000010101010011;
            15'd21973: log10_cal = 16'b0000010101010011;
            15'd21974: log10_cal = 16'b0000010101010011;
            15'd21975: log10_cal = 16'b0000010101010011;
            15'd21976: log10_cal = 16'b0000010101010011;
            15'd21977: log10_cal = 16'b0000010101010011;
            15'd21978: log10_cal = 16'b0000010101010011;
            15'd21979: log10_cal = 16'b0000010101010011;
            15'd21980: log10_cal = 16'b0000010101010011;
            15'd21981: log10_cal = 16'b0000010101010011;
            15'd21982: log10_cal = 16'b0000010101010011;
            15'd21983: log10_cal = 16'b0000010101010011;
            15'd21984: log10_cal = 16'b0000010101010011;
            15'd21985: log10_cal = 16'b0000010101010011;
            15'd21986: log10_cal = 16'b0000010101010011;
            15'd21987: log10_cal = 16'b0000010101010011;
            15'd21988: log10_cal = 16'b0000010101010011;
            15'd21989: log10_cal = 16'b0000010101010011;
            15'd21990: log10_cal = 16'b0000010101010011;
            15'd21991: log10_cal = 16'b0000010101010011;
            15'd21992: log10_cal = 16'b0000010101010011;
            15'd21993: log10_cal = 16'b0000010101010011;
            15'd21994: log10_cal = 16'b0000010101010011;
            15'd21995: log10_cal = 16'b0000010101010011;
            15'd21996: log10_cal = 16'b0000010101010100;
            15'd21997: log10_cal = 16'b0000010101010100;
            15'd21998: log10_cal = 16'b0000010101010100;
            15'd21999: log10_cal = 16'b0000010101010100;
            15'd22000: log10_cal = 16'b0000010101010100;
            15'd22001: log10_cal = 16'b0000010101010100;
            15'd22002: log10_cal = 16'b0000010101010100;
            15'd22003: log10_cal = 16'b0000010101010100;
            15'd22004: log10_cal = 16'b0000010101010100;
            15'd22005: log10_cal = 16'b0000010101010100;
            15'd22006: log10_cal = 16'b0000010101010100;
            15'd22007: log10_cal = 16'b0000010101010100;
            15'd22008: log10_cal = 16'b0000010101010100;
            15'd22009: log10_cal = 16'b0000010101010100;
            15'd22010: log10_cal = 16'b0000010101010100;
            15'd22011: log10_cal = 16'b0000010101010100;
            15'd22012: log10_cal = 16'b0000010101010100;
            15'd22013: log10_cal = 16'b0000010101010100;
            15'd22014: log10_cal = 16'b0000010101010100;
            15'd22015: log10_cal = 16'b0000010101010100;
            15'd22016: log10_cal = 16'b0000010101010100;
            15'd22017: log10_cal = 16'b0000010101010100;
            15'd22018: log10_cal = 16'b0000010101010100;
            15'd22019: log10_cal = 16'b0000010101010100;
            15'd22020: log10_cal = 16'b0000010101010100;
            15'd22021: log10_cal = 16'b0000010101010100;
            15'd22022: log10_cal = 16'b0000010101010100;
            15'd22023: log10_cal = 16'b0000010101010100;
            15'd22024: log10_cal = 16'b0000010101010100;
            15'd22025: log10_cal = 16'b0000010101010100;
            15'd22026: log10_cal = 16'b0000010101010100;
            15'd22027: log10_cal = 16'b0000010101010100;
            15'd22028: log10_cal = 16'b0000010101010100;
            15'd22029: log10_cal = 16'b0000010101010100;
            15'd22030: log10_cal = 16'b0000010101010100;
            15'd22031: log10_cal = 16'b0000010101010100;
            15'd22032: log10_cal = 16'b0000010101010100;
            15'd22033: log10_cal = 16'b0000010101010100;
            15'd22034: log10_cal = 16'b0000010101010100;
            15'd22035: log10_cal = 16'b0000010101010100;
            15'd22036: log10_cal = 16'b0000010101010100;
            15'd22037: log10_cal = 16'b0000010101010100;
            15'd22038: log10_cal = 16'b0000010101010100;
            15'd22039: log10_cal = 16'b0000010101010100;
            15'd22040: log10_cal = 16'b0000010101010100;
            15'd22041: log10_cal = 16'b0000010101010100;
            15'd22042: log10_cal = 16'b0000010101010100;
            15'd22043: log10_cal = 16'b0000010101010100;
            15'd22044: log10_cal = 16'b0000010101010100;
            15'd22045: log10_cal = 16'b0000010101010101;
            15'd22046: log10_cal = 16'b0000010101010101;
            15'd22047: log10_cal = 16'b0000010101010101;
            15'd22048: log10_cal = 16'b0000010101010101;
            15'd22049: log10_cal = 16'b0000010101010101;
            15'd22050: log10_cal = 16'b0000010101010101;
            15'd22051: log10_cal = 16'b0000010101010101;
            15'd22052: log10_cal = 16'b0000010101010101;
            15'd22053: log10_cal = 16'b0000010101010101;
            15'd22054: log10_cal = 16'b0000010101010101;
            15'd22055: log10_cal = 16'b0000010101010101;
            15'd22056: log10_cal = 16'b0000010101010101;
            15'd22057: log10_cal = 16'b0000010101010101;
            15'd22058: log10_cal = 16'b0000010101010101;
            15'd22059: log10_cal = 16'b0000010101010101;
            15'd22060: log10_cal = 16'b0000010101010101;
            15'd22061: log10_cal = 16'b0000010101010101;
            15'd22062: log10_cal = 16'b0000010101010101;
            15'd22063: log10_cal = 16'b0000010101010101;
            15'd22064: log10_cal = 16'b0000010101010101;
            15'd22065: log10_cal = 16'b0000010101010101;
            15'd22066: log10_cal = 16'b0000010101010101;
            15'd22067: log10_cal = 16'b0000010101010101;
            15'd22068: log10_cal = 16'b0000010101010101;
            15'd22069: log10_cal = 16'b0000010101010101;
            15'd22070: log10_cal = 16'b0000010101010101;
            15'd22071: log10_cal = 16'b0000010101010101;
            15'd22072: log10_cal = 16'b0000010101010101;
            15'd22073: log10_cal = 16'b0000010101010101;
            15'd22074: log10_cal = 16'b0000010101010101;
            15'd22075: log10_cal = 16'b0000010101010101;
            15'd22076: log10_cal = 16'b0000010101010101;
            15'd22077: log10_cal = 16'b0000010101010101;
            15'd22078: log10_cal = 16'b0000010101010101;
            15'd22079: log10_cal = 16'b0000010101010101;
            15'd22080: log10_cal = 16'b0000010101010101;
            15'd22081: log10_cal = 16'b0000010101010101;
            15'd22082: log10_cal = 16'b0000010101010101;
            15'd22083: log10_cal = 16'b0000010101010101;
            15'd22084: log10_cal = 16'b0000010101010101;
            15'd22085: log10_cal = 16'b0000010101010101;
            15'd22086: log10_cal = 16'b0000010101010101;
            15'd22087: log10_cal = 16'b0000010101010101;
            15'd22088: log10_cal = 16'b0000010101010101;
            15'd22089: log10_cal = 16'b0000010101010101;
            15'd22090: log10_cal = 16'b0000010101010101;
            15'd22091: log10_cal = 16'b0000010101010101;
            15'd22092: log10_cal = 16'b0000010101010101;
            15'd22093: log10_cal = 16'b0000010101010101;
            15'd22094: log10_cal = 16'b0000010101010101;
            15'd22095: log10_cal = 16'b0000010101010110;
            15'd22096: log10_cal = 16'b0000010101010110;
            15'd22097: log10_cal = 16'b0000010101010110;
            15'd22098: log10_cal = 16'b0000010101010110;
            15'd22099: log10_cal = 16'b0000010101010110;
            15'd22100: log10_cal = 16'b0000010101010110;
            15'd22101: log10_cal = 16'b0000010101010110;
            15'd22102: log10_cal = 16'b0000010101010110;
            15'd22103: log10_cal = 16'b0000010101010110;
            15'd22104: log10_cal = 16'b0000010101010110;
            15'd22105: log10_cal = 16'b0000010101010110;
            15'd22106: log10_cal = 16'b0000010101010110;
            15'd22107: log10_cal = 16'b0000010101010110;
            15'd22108: log10_cal = 16'b0000010101010110;
            15'd22109: log10_cal = 16'b0000010101010110;
            15'd22110: log10_cal = 16'b0000010101010110;
            15'd22111: log10_cal = 16'b0000010101010110;
            15'd22112: log10_cal = 16'b0000010101010110;
            15'd22113: log10_cal = 16'b0000010101010110;
            15'd22114: log10_cal = 16'b0000010101010110;
            15'd22115: log10_cal = 16'b0000010101010110;
            15'd22116: log10_cal = 16'b0000010101010110;
            15'd22117: log10_cal = 16'b0000010101010110;
            15'd22118: log10_cal = 16'b0000010101010110;
            15'd22119: log10_cal = 16'b0000010101010110;
            15'd22120: log10_cal = 16'b0000010101010110;
            15'd22121: log10_cal = 16'b0000010101010110;
            15'd22122: log10_cal = 16'b0000010101010110;
            15'd22123: log10_cal = 16'b0000010101010110;
            15'd22124: log10_cal = 16'b0000010101010110;
            15'd22125: log10_cal = 16'b0000010101010110;
            15'd22126: log10_cal = 16'b0000010101010110;
            15'd22127: log10_cal = 16'b0000010101010110;
            15'd22128: log10_cal = 16'b0000010101010110;
            15'd22129: log10_cal = 16'b0000010101010110;
            15'd22130: log10_cal = 16'b0000010101010110;
            15'd22131: log10_cal = 16'b0000010101010110;
            15'd22132: log10_cal = 16'b0000010101010110;
            15'd22133: log10_cal = 16'b0000010101010110;
            15'd22134: log10_cal = 16'b0000010101010110;
            15'd22135: log10_cal = 16'b0000010101010110;
            15'd22136: log10_cal = 16'b0000010101010110;
            15'd22137: log10_cal = 16'b0000010101010110;
            15'd22138: log10_cal = 16'b0000010101010110;
            15'd22139: log10_cal = 16'b0000010101010110;
            15'd22140: log10_cal = 16'b0000010101010110;
            15'd22141: log10_cal = 16'b0000010101010110;
            15'd22142: log10_cal = 16'b0000010101010110;
            15'd22143: log10_cal = 16'b0000010101010110;
            15'd22144: log10_cal = 16'b0000010101010110;
            15'd22145: log10_cal = 16'b0000010101010111;
            15'd22146: log10_cal = 16'b0000010101010111;
            15'd22147: log10_cal = 16'b0000010101010111;
            15'd22148: log10_cal = 16'b0000010101010111;
            15'd22149: log10_cal = 16'b0000010101010111;
            15'd22150: log10_cal = 16'b0000010101010111;
            15'd22151: log10_cal = 16'b0000010101010111;
            15'd22152: log10_cal = 16'b0000010101010111;
            15'd22153: log10_cal = 16'b0000010101010111;
            15'd22154: log10_cal = 16'b0000010101010111;
            15'd22155: log10_cal = 16'b0000010101010111;
            15'd22156: log10_cal = 16'b0000010101010111;
            15'd22157: log10_cal = 16'b0000010101010111;
            15'd22158: log10_cal = 16'b0000010101010111;
            15'd22159: log10_cal = 16'b0000010101010111;
            15'd22160: log10_cal = 16'b0000010101010111;
            15'd22161: log10_cal = 16'b0000010101010111;
            15'd22162: log10_cal = 16'b0000010101010111;
            15'd22163: log10_cal = 16'b0000010101010111;
            15'd22164: log10_cal = 16'b0000010101010111;
            15'd22165: log10_cal = 16'b0000010101010111;
            15'd22166: log10_cal = 16'b0000010101010111;
            15'd22167: log10_cal = 16'b0000010101010111;
            15'd22168: log10_cal = 16'b0000010101010111;
            15'd22169: log10_cal = 16'b0000010101010111;
            15'd22170: log10_cal = 16'b0000010101010111;
            15'd22171: log10_cal = 16'b0000010101010111;
            15'd22172: log10_cal = 16'b0000010101010111;
            15'd22173: log10_cal = 16'b0000010101010111;
            15'd22174: log10_cal = 16'b0000010101010111;
            15'd22175: log10_cal = 16'b0000010101010111;
            15'd22176: log10_cal = 16'b0000010101010111;
            15'd22177: log10_cal = 16'b0000010101010111;
            15'd22178: log10_cal = 16'b0000010101010111;
            15'd22179: log10_cal = 16'b0000010101010111;
            15'd22180: log10_cal = 16'b0000010101010111;
            15'd22181: log10_cal = 16'b0000010101010111;
            15'd22182: log10_cal = 16'b0000010101010111;
            15'd22183: log10_cal = 16'b0000010101010111;
            15'd22184: log10_cal = 16'b0000010101010111;
            15'd22185: log10_cal = 16'b0000010101010111;
            15'd22186: log10_cal = 16'b0000010101010111;
            15'd22187: log10_cal = 16'b0000010101010111;
            15'd22188: log10_cal = 16'b0000010101010111;
            15'd22189: log10_cal = 16'b0000010101010111;
            15'd22190: log10_cal = 16'b0000010101010111;
            15'd22191: log10_cal = 16'b0000010101010111;
            15'd22192: log10_cal = 16'b0000010101010111;
            15'd22193: log10_cal = 16'b0000010101010111;
            15'd22194: log10_cal = 16'b0000010101010111;
            15'd22195: log10_cal = 16'b0000010101011000;
            15'd22196: log10_cal = 16'b0000010101011000;
            15'd22197: log10_cal = 16'b0000010101011000;
            15'd22198: log10_cal = 16'b0000010101011000;
            15'd22199: log10_cal = 16'b0000010101011000;
            15'd22200: log10_cal = 16'b0000010101011000;
            15'd22201: log10_cal = 16'b0000010101011000;
            15'd22202: log10_cal = 16'b0000010101011000;
            15'd22203: log10_cal = 16'b0000010101011000;
            15'd22204: log10_cal = 16'b0000010101011000;
            15'd22205: log10_cal = 16'b0000010101011000;
            15'd22206: log10_cal = 16'b0000010101011000;
            15'd22207: log10_cal = 16'b0000010101011000;
            15'd22208: log10_cal = 16'b0000010101011000;
            15'd22209: log10_cal = 16'b0000010101011000;
            15'd22210: log10_cal = 16'b0000010101011000;
            15'd22211: log10_cal = 16'b0000010101011000;
            15'd22212: log10_cal = 16'b0000010101011000;
            15'd22213: log10_cal = 16'b0000010101011000;
            15'd22214: log10_cal = 16'b0000010101011000;
            15'd22215: log10_cal = 16'b0000010101011000;
            15'd22216: log10_cal = 16'b0000010101011000;
            15'd22217: log10_cal = 16'b0000010101011000;
            15'd22218: log10_cal = 16'b0000010101011000;
            15'd22219: log10_cal = 16'b0000010101011000;
            15'd22220: log10_cal = 16'b0000010101011000;
            15'd22221: log10_cal = 16'b0000010101011000;
            15'd22222: log10_cal = 16'b0000010101011000;
            15'd22223: log10_cal = 16'b0000010101011000;
            15'd22224: log10_cal = 16'b0000010101011000;
            15'd22225: log10_cal = 16'b0000010101011000;
            15'd22226: log10_cal = 16'b0000010101011000;
            15'd22227: log10_cal = 16'b0000010101011000;
            15'd22228: log10_cal = 16'b0000010101011000;
            15'd22229: log10_cal = 16'b0000010101011000;
            15'd22230: log10_cal = 16'b0000010101011000;
            15'd22231: log10_cal = 16'b0000010101011000;
            15'd22232: log10_cal = 16'b0000010101011000;
            15'd22233: log10_cal = 16'b0000010101011000;
            15'd22234: log10_cal = 16'b0000010101011000;
            15'd22235: log10_cal = 16'b0000010101011000;
            15'd22236: log10_cal = 16'b0000010101011000;
            15'd22237: log10_cal = 16'b0000010101011000;
            15'd22238: log10_cal = 16'b0000010101011000;
            15'd22239: log10_cal = 16'b0000010101011000;
            15'd22240: log10_cal = 16'b0000010101011000;
            15'd22241: log10_cal = 16'b0000010101011000;
            15'd22242: log10_cal = 16'b0000010101011000;
            15'd22243: log10_cal = 16'b0000010101011000;
            15'd22244: log10_cal = 16'b0000010101011000;
            15'd22245: log10_cal = 16'b0000010101011001;
            15'd22246: log10_cal = 16'b0000010101011001;
            15'd22247: log10_cal = 16'b0000010101011001;
            15'd22248: log10_cal = 16'b0000010101011001;
            15'd22249: log10_cal = 16'b0000010101011001;
            15'd22250: log10_cal = 16'b0000010101011001;
            15'd22251: log10_cal = 16'b0000010101011001;
            15'd22252: log10_cal = 16'b0000010101011001;
            15'd22253: log10_cal = 16'b0000010101011001;
            15'd22254: log10_cal = 16'b0000010101011001;
            15'd22255: log10_cal = 16'b0000010101011001;
            15'd22256: log10_cal = 16'b0000010101011001;
            15'd22257: log10_cal = 16'b0000010101011001;
            15'd22258: log10_cal = 16'b0000010101011001;
            15'd22259: log10_cal = 16'b0000010101011001;
            15'd22260: log10_cal = 16'b0000010101011001;
            15'd22261: log10_cal = 16'b0000010101011001;
            15'd22262: log10_cal = 16'b0000010101011001;
            15'd22263: log10_cal = 16'b0000010101011001;
            15'd22264: log10_cal = 16'b0000010101011001;
            15'd22265: log10_cal = 16'b0000010101011001;
            15'd22266: log10_cal = 16'b0000010101011001;
            15'd22267: log10_cal = 16'b0000010101011001;
            15'd22268: log10_cal = 16'b0000010101011001;
            15'd22269: log10_cal = 16'b0000010101011001;
            15'd22270: log10_cal = 16'b0000010101011001;
            15'd22271: log10_cal = 16'b0000010101011001;
            15'd22272: log10_cal = 16'b0000010101011001;
            15'd22273: log10_cal = 16'b0000010101011001;
            15'd22274: log10_cal = 16'b0000010101011001;
            15'd22275: log10_cal = 16'b0000010101011001;
            15'd22276: log10_cal = 16'b0000010101011001;
            15'd22277: log10_cal = 16'b0000010101011001;
            15'd22278: log10_cal = 16'b0000010101011001;
            15'd22279: log10_cal = 16'b0000010101011001;
            15'd22280: log10_cal = 16'b0000010101011001;
            15'd22281: log10_cal = 16'b0000010101011001;
            15'd22282: log10_cal = 16'b0000010101011001;
            15'd22283: log10_cal = 16'b0000010101011001;
            15'd22284: log10_cal = 16'b0000010101011001;
            15'd22285: log10_cal = 16'b0000010101011001;
            15'd22286: log10_cal = 16'b0000010101011001;
            15'd22287: log10_cal = 16'b0000010101011001;
            15'd22288: log10_cal = 16'b0000010101011001;
            15'd22289: log10_cal = 16'b0000010101011001;
            15'd22290: log10_cal = 16'b0000010101011001;
            15'd22291: log10_cal = 16'b0000010101011001;
            15'd22292: log10_cal = 16'b0000010101011001;
            15'd22293: log10_cal = 16'b0000010101011001;
            15'd22294: log10_cal = 16'b0000010101011001;
            15'd22295: log10_cal = 16'b0000010101011010;
            15'd22296: log10_cal = 16'b0000010101011010;
            15'd22297: log10_cal = 16'b0000010101011010;
            15'd22298: log10_cal = 16'b0000010101011010;
            15'd22299: log10_cal = 16'b0000010101011010;
            15'd22300: log10_cal = 16'b0000010101011010;
            15'd22301: log10_cal = 16'b0000010101011010;
            15'd22302: log10_cal = 16'b0000010101011010;
            15'd22303: log10_cal = 16'b0000010101011010;
            15'd22304: log10_cal = 16'b0000010101011010;
            15'd22305: log10_cal = 16'b0000010101011010;
            15'd22306: log10_cal = 16'b0000010101011010;
            15'd22307: log10_cal = 16'b0000010101011010;
            15'd22308: log10_cal = 16'b0000010101011010;
            15'd22309: log10_cal = 16'b0000010101011010;
            15'd22310: log10_cal = 16'b0000010101011010;
            15'd22311: log10_cal = 16'b0000010101011010;
            15'd22312: log10_cal = 16'b0000010101011010;
            15'd22313: log10_cal = 16'b0000010101011010;
            15'd22314: log10_cal = 16'b0000010101011010;
            15'd22315: log10_cal = 16'b0000010101011010;
            15'd22316: log10_cal = 16'b0000010101011010;
            15'd22317: log10_cal = 16'b0000010101011010;
            15'd22318: log10_cal = 16'b0000010101011010;
            15'd22319: log10_cal = 16'b0000010101011010;
            15'd22320: log10_cal = 16'b0000010101011010;
            15'd22321: log10_cal = 16'b0000010101011010;
            15'd22322: log10_cal = 16'b0000010101011010;
            15'd22323: log10_cal = 16'b0000010101011010;
            15'd22324: log10_cal = 16'b0000010101011010;
            15'd22325: log10_cal = 16'b0000010101011010;
            15'd22326: log10_cal = 16'b0000010101011010;
            15'd22327: log10_cal = 16'b0000010101011010;
            15'd22328: log10_cal = 16'b0000010101011010;
            15'd22329: log10_cal = 16'b0000010101011010;
            15'd22330: log10_cal = 16'b0000010101011010;
            15'd22331: log10_cal = 16'b0000010101011010;
            15'd22332: log10_cal = 16'b0000010101011010;
            15'd22333: log10_cal = 16'b0000010101011010;
            15'd22334: log10_cal = 16'b0000010101011010;
            15'd22335: log10_cal = 16'b0000010101011010;
            15'd22336: log10_cal = 16'b0000010101011010;
            15'd22337: log10_cal = 16'b0000010101011010;
            15'd22338: log10_cal = 16'b0000010101011010;
            15'd22339: log10_cal = 16'b0000010101011010;
            15'd22340: log10_cal = 16'b0000010101011010;
            15'd22341: log10_cal = 16'b0000010101011010;
            15'd22342: log10_cal = 16'b0000010101011010;
            15'd22343: log10_cal = 16'b0000010101011010;
            15'd22344: log10_cal = 16'b0000010101011010;
            15'd22345: log10_cal = 16'b0000010101011011;
            15'd22346: log10_cal = 16'b0000010101011011;
            15'd22347: log10_cal = 16'b0000010101011011;
            15'd22348: log10_cal = 16'b0000010101011011;
            15'd22349: log10_cal = 16'b0000010101011011;
            15'd22350: log10_cal = 16'b0000010101011011;
            15'd22351: log10_cal = 16'b0000010101011011;
            15'd22352: log10_cal = 16'b0000010101011011;
            15'd22353: log10_cal = 16'b0000010101011011;
            15'd22354: log10_cal = 16'b0000010101011011;
            15'd22355: log10_cal = 16'b0000010101011011;
            15'd22356: log10_cal = 16'b0000010101011011;
            15'd22357: log10_cal = 16'b0000010101011011;
            15'd22358: log10_cal = 16'b0000010101011011;
            15'd22359: log10_cal = 16'b0000010101011011;
            15'd22360: log10_cal = 16'b0000010101011011;
            15'd22361: log10_cal = 16'b0000010101011011;
            15'd22362: log10_cal = 16'b0000010101011011;
            15'd22363: log10_cal = 16'b0000010101011011;
            15'd22364: log10_cal = 16'b0000010101011011;
            15'd22365: log10_cal = 16'b0000010101011011;
            15'd22366: log10_cal = 16'b0000010101011011;
            15'd22367: log10_cal = 16'b0000010101011011;
            15'd22368: log10_cal = 16'b0000010101011011;
            15'd22369: log10_cal = 16'b0000010101011011;
            15'd22370: log10_cal = 16'b0000010101011011;
            15'd22371: log10_cal = 16'b0000010101011011;
            15'd22372: log10_cal = 16'b0000010101011011;
            15'd22373: log10_cal = 16'b0000010101011011;
            15'd22374: log10_cal = 16'b0000010101011011;
            15'd22375: log10_cal = 16'b0000010101011011;
            15'd22376: log10_cal = 16'b0000010101011011;
            15'd22377: log10_cal = 16'b0000010101011011;
            15'd22378: log10_cal = 16'b0000010101011011;
            15'd22379: log10_cal = 16'b0000010101011011;
            15'd22380: log10_cal = 16'b0000010101011011;
            15'd22381: log10_cal = 16'b0000010101011011;
            15'd22382: log10_cal = 16'b0000010101011011;
            15'd22383: log10_cal = 16'b0000010101011011;
            15'd22384: log10_cal = 16'b0000010101011011;
            15'd22385: log10_cal = 16'b0000010101011011;
            15'd22386: log10_cal = 16'b0000010101011011;
            15'd22387: log10_cal = 16'b0000010101011011;
            15'd22388: log10_cal = 16'b0000010101011011;
            15'd22389: log10_cal = 16'b0000010101011011;
            15'd22390: log10_cal = 16'b0000010101011011;
            15'd22391: log10_cal = 16'b0000010101011011;
            15'd22392: log10_cal = 16'b0000010101011011;
            15'd22393: log10_cal = 16'b0000010101011011;
            15'd22394: log10_cal = 16'b0000010101011011;
            15'd22395: log10_cal = 16'b0000010101011100;
            15'd22396: log10_cal = 16'b0000010101011100;
            15'd22397: log10_cal = 16'b0000010101011100;
            15'd22398: log10_cal = 16'b0000010101011100;
            15'd22399: log10_cal = 16'b0000010101011100;
            15'd22400: log10_cal = 16'b0000010101011100;
            15'd22401: log10_cal = 16'b0000010101011100;
            15'd22402: log10_cal = 16'b0000010101011100;
            15'd22403: log10_cal = 16'b0000010101011100;
            15'd22404: log10_cal = 16'b0000010101011100;
            15'd22405: log10_cal = 16'b0000010101011100;
            15'd22406: log10_cal = 16'b0000010101011100;
            15'd22407: log10_cal = 16'b0000010101011100;
            15'd22408: log10_cal = 16'b0000010101011100;
            15'd22409: log10_cal = 16'b0000010101011100;
            15'd22410: log10_cal = 16'b0000010101011100;
            15'd22411: log10_cal = 16'b0000010101011100;
            15'd22412: log10_cal = 16'b0000010101011100;
            15'd22413: log10_cal = 16'b0000010101011100;
            15'd22414: log10_cal = 16'b0000010101011100;
            15'd22415: log10_cal = 16'b0000010101011100;
            15'd22416: log10_cal = 16'b0000010101011100;
            15'd22417: log10_cal = 16'b0000010101011100;
            15'd22418: log10_cal = 16'b0000010101011100;
            15'd22419: log10_cal = 16'b0000010101011100;
            15'd22420: log10_cal = 16'b0000010101011100;
            15'd22421: log10_cal = 16'b0000010101011100;
            15'd22422: log10_cal = 16'b0000010101011100;
            15'd22423: log10_cal = 16'b0000010101011100;
            15'd22424: log10_cal = 16'b0000010101011100;
            15'd22425: log10_cal = 16'b0000010101011100;
            15'd22426: log10_cal = 16'b0000010101011100;
            15'd22427: log10_cal = 16'b0000010101011100;
            15'd22428: log10_cal = 16'b0000010101011100;
            15'd22429: log10_cal = 16'b0000010101011100;
            15'd22430: log10_cal = 16'b0000010101011100;
            15'd22431: log10_cal = 16'b0000010101011100;
            15'd22432: log10_cal = 16'b0000010101011100;
            15'd22433: log10_cal = 16'b0000010101011100;
            15'd22434: log10_cal = 16'b0000010101011100;
            15'd22435: log10_cal = 16'b0000010101011100;
            15'd22436: log10_cal = 16'b0000010101011100;
            15'd22437: log10_cal = 16'b0000010101011100;
            15'd22438: log10_cal = 16'b0000010101011100;
            15'd22439: log10_cal = 16'b0000010101011100;
            15'd22440: log10_cal = 16'b0000010101011100;
            15'd22441: log10_cal = 16'b0000010101011100;
            15'd22442: log10_cal = 16'b0000010101011100;
            15'd22443: log10_cal = 16'b0000010101011100;
            15'd22444: log10_cal = 16'b0000010101011100;
            15'd22445: log10_cal = 16'b0000010101011100;
            15'd22446: log10_cal = 16'b0000010101011101;
            15'd22447: log10_cal = 16'b0000010101011101;
            15'd22448: log10_cal = 16'b0000010101011101;
            15'd22449: log10_cal = 16'b0000010101011101;
            15'd22450: log10_cal = 16'b0000010101011101;
            15'd22451: log10_cal = 16'b0000010101011101;
            15'd22452: log10_cal = 16'b0000010101011101;
            15'd22453: log10_cal = 16'b0000010101011101;
            15'd22454: log10_cal = 16'b0000010101011101;
            15'd22455: log10_cal = 16'b0000010101011101;
            15'd22456: log10_cal = 16'b0000010101011101;
            15'd22457: log10_cal = 16'b0000010101011101;
            15'd22458: log10_cal = 16'b0000010101011101;
            15'd22459: log10_cal = 16'b0000010101011101;
            15'd22460: log10_cal = 16'b0000010101011101;
            15'd22461: log10_cal = 16'b0000010101011101;
            15'd22462: log10_cal = 16'b0000010101011101;
            15'd22463: log10_cal = 16'b0000010101011101;
            15'd22464: log10_cal = 16'b0000010101011101;
            15'd22465: log10_cal = 16'b0000010101011101;
            15'd22466: log10_cal = 16'b0000010101011101;
            15'd22467: log10_cal = 16'b0000010101011101;
            15'd22468: log10_cal = 16'b0000010101011101;
            15'd22469: log10_cal = 16'b0000010101011101;
            15'd22470: log10_cal = 16'b0000010101011101;
            15'd22471: log10_cal = 16'b0000010101011101;
            15'd22472: log10_cal = 16'b0000010101011101;
            15'd22473: log10_cal = 16'b0000010101011101;
            15'd22474: log10_cal = 16'b0000010101011101;
            15'd22475: log10_cal = 16'b0000010101011101;
            15'd22476: log10_cal = 16'b0000010101011101;
            15'd22477: log10_cal = 16'b0000010101011101;
            15'd22478: log10_cal = 16'b0000010101011101;
            15'd22479: log10_cal = 16'b0000010101011101;
            15'd22480: log10_cal = 16'b0000010101011101;
            15'd22481: log10_cal = 16'b0000010101011101;
            15'd22482: log10_cal = 16'b0000010101011101;
            15'd22483: log10_cal = 16'b0000010101011101;
            15'd22484: log10_cal = 16'b0000010101011101;
            15'd22485: log10_cal = 16'b0000010101011101;
            15'd22486: log10_cal = 16'b0000010101011101;
            15'd22487: log10_cal = 16'b0000010101011101;
            15'd22488: log10_cal = 16'b0000010101011101;
            15'd22489: log10_cal = 16'b0000010101011101;
            15'd22490: log10_cal = 16'b0000010101011101;
            15'd22491: log10_cal = 16'b0000010101011101;
            15'd22492: log10_cal = 16'b0000010101011101;
            15'd22493: log10_cal = 16'b0000010101011101;
            15'd22494: log10_cal = 16'b0000010101011101;
            15'd22495: log10_cal = 16'b0000010101011101;
            15'd22496: log10_cal = 16'b0000010101011110;
            15'd22497: log10_cal = 16'b0000010101011110;
            15'd22498: log10_cal = 16'b0000010101011110;
            15'd22499: log10_cal = 16'b0000010101011110;
            15'd22500: log10_cal = 16'b0000010101011110;
            15'd22501: log10_cal = 16'b0000010101011110;
            15'd22502: log10_cal = 16'b0000010101011110;
            15'd22503: log10_cal = 16'b0000010101011110;
            15'd22504: log10_cal = 16'b0000010101011110;
            15'd22505: log10_cal = 16'b0000010101011110;
            15'd22506: log10_cal = 16'b0000010101011110;
            15'd22507: log10_cal = 16'b0000010101011110;
            15'd22508: log10_cal = 16'b0000010101011110;
            15'd22509: log10_cal = 16'b0000010101011110;
            15'd22510: log10_cal = 16'b0000010101011110;
            15'd22511: log10_cal = 16'b0000010101011110;
            15'd22512: log10_cal = 16'b0000010101011110;
            15'd22513: log10_cal = 16'b0000010101011110;
            15'd22514: log10_cal = 16'b0000010101011110;
            15'd22515: log10_cal = 16'b0000010101011110;
            15'd22516: log10_cal = 16'b0000010101011110;
            15'd22517: log10_cal = 16'b0000010101011110;
            15'd22518: log10_cal = 16'b0000010101011110;
            15'd22519: log10_cal = 16'b0000010101011110;
            15'd22520: log10_cal = 16'b0000010101011110;
            15'd22521: log10_cal = 16'b0000010101011110;
            15'd22522: log10_cal = 16'b0000010101011110;
            15'd22523: log10_cal = 16'b0000010101011110;
            15'd22524: log10_cal = 16'b0000010101011110;
            15'd22525: log10_cal = 16'b0000010101011110;
            15'd22526: log10_cal = 16'b0000010101011110;
            15'd22527: log10_cal = 16'b0000010101011110;
            15'd22528: log10_cal = 16'b0000010101011110;
            15'd22529: log10_cal = 16'b0000010101011110;
            15'd22530: log10_cal = 16'b0000010101011110;
            15'd22531: log10_cal = 16'b0000010101011110;
            15'd22532: log10_cal = 16'b0000010101011110;
            15'd22533: log10_cal = 16'b0000010101011110;
            15'd22534: log10_cal = 16'b0000010101011110;
            15'd22535: log10_cal = 16'b0000010101011110;
            15'd22536: log10_cal = 16'b0000010101011110;
            15'd22537: log10_cal = 16'b0000010101011110;
            15'd22538: log10_cal = 16'b0000010101011110;
            15'd22539: log10_cal = 16'b0000010101011110;
            15'd22540: log10_cal = 16'b0000010101011110;
            15'd22541: log10_cal = 16'b0000010101011110;
            15'd22542: log10_cal = 16'b0000010101011110;
            15'd22543: log10_cal = 16'b0000010101011110;
            15'd22544: log10_cal = 16'b0000010101011110;
            15'd22545: log10_cal = 16'b0000010101011110;
            15'd22546: log10_cal = 16'b0000010101011110;
            15'd22547: log10_cal = 16'b0000010101011111;
            15'd22548: log10_cal = 16'b0000010101011111;
            15'd22549: log10_cal = 16'b0000010101011111;
            15'd22550: log10_cal = 16'b0000010101011111;
            15'd22551: log10_cal = 16'b0000010101011111;
            15'd22552: log10_cal = 16'b0000010101011111;
            15'd22553: log10_cal = 16'b0000010101011111;
            15'd22554: log10_cal = 16'b0000010101011111;
            15'd22555: log10_cal = 16'b0000010101011111;
            15'd22556: log10_cal = 16'b0000010101011111;
            15'd22557: log10_cal = 16'b0000010101011111;
            15'd22558: log10_cal = 16'b0000010101011111;
            15'd22559: log10_cal = 16'b0000010101011111;
            15'd22560: log10_cal = 16'b0000010101011111;
            15'd22561: log10_cal = 16'b0000010101011111;
            15'd22562: log10_cal = 16'b0000010101011111;
            15'd22563: log10_cal = 16'b0000010101011111;
            15'd22564: log10_cal = 16'b0000010101011111;
            15'd22565: log10_cal = 16'b0000010101011111;
            15'd22566: log10_cal = 16'b0000010101011111;
            15'd22567: log10_cal = 16'b0000010101011111;
            15'd22568: log10_cal = 16'b0000010101011111;
            15'd22569: log10_cal = 16'b0000010101011111;
            15'd22570: log10_cal = 16'b0000010101011111;
            15'd22571: log10_cal = 16'b0000010101011111;
            15'd22572: log10_cal = 16'b0000010101011111;
            15'd22573: log10_cal = 16'b0000010101011111;
            15'd22574: log10_cal = 16'b0000010101011111;
            15'd22575: log10_cal = 16'b0000010101011111;
            15'd22576: log10_cal = 16'b0000010101011111;
            15'd22577: log10_cal = 16'b0000010101011111;
            15'd22578: log10_cal = 16'b0000010101011111;
            15'd22579: log10_cal = 16'b0000010101011111;
            15'd22580: log10_cal = 16'b0000010101011111;
            15'd22581: log10_cal = 16'b0000010101011111;
            15'd22582: log10_cal = 16'b0000010101011111;
            15'd22583: log10_cal = 16'b0000010101011111;
            15'd22584: log10_cal = 16'b0000010101011111;
            15'd22585: log10_cal = 16'b0000010101011111;
            15'd22586: log10_cal = 16'b0000010101011111;
            15'd22587: log10_cal = 16'b0000010101011111;
            15'd22588: log10_cal = 16'b0000010101011111;
            15'd22589: log10_cal = 16'b0000010101011111;
            15'd22590: log10_cal = 16'b0000010101011111;
            15'd22591: log10_cal = 16'b0000010101011111;
            15'd22592: log10_cal = 16'b0000010101011111;
            15'd22593: log10_cal = 16'b0000010101011111;
            15'd22594: log10_cal = 16'b0000010101011111;
            15'd22595: log10_cal = 16'b0000010101011111;
            15'd22596: log10_cal = 16'b0000010101011111;
            15'd22597: log10_cal = 16'b0000010101100000;
            15'd22598: log10_cal = 16'b0000010101100000;
            15'd22599: log10_cal = 16'b0000010101100000;
            15'd22600: log10_cal = 16'b0000010101100000;
            15'd22601: log10_cal = 16'b0000010101100000;
            15'd22602: log10_cal = 16'b0000010101100000;
            15'd22603: log10_cal = 16'b0000010101100000;
            15'd22604: log10_cal = 16'b0000010101100000;
            15'd22605: log10_cal = 16'b0000010101100000;
            15'd22606: log10_cal = 16'b0000010101100000;
            15'd22607: log10_cal = 16'b0000010101100000;
            15'd22608: log10_cal = 16'b0000010101100000;
            15'd22609: log10_cal = 16'b0000010101100000;
            15'd22610: log10_cal = 16'b0000010101100000;
            15'd22611: log10_cal = 16'b0000010101100000;
            15'd22612: log10_cal = 16'b0000010101100000;
            15'd22613: log10_cal = 16'b0000010101100000;
            15'd22614: log10_cal = 16'b0000010101100000;
            15'd22615: log10_cal = 16'b0000010101100000;
            15'd22616: log10_cal = 16'b0000010101100000;
            15'd22617: log10_cal = 16'b0000010101100000;
            15'd22618: log10_cal = 16'b0000010101100000;
            15'd22619: log10_cal = 16'b0000010101100000;
            15'd22620: log10_cal = 16'b0000010101100000;
            15'd22621: log10_cal = 16'b0000010101100000;
            15'd22622: log10_cal = 16'b0000010101100000;
            15'd22623: log10_cal = 16'b0000010101100000;
            15'd22624: log10_cal = 16'b0000010101100000;
            15'd22625: log10_cal = 16'b0000010101100000;
            15'd22626: log10_cal = 16'b0000010101100000;
            15'd22627: log10_cal = 16'b0000010101100000;
            15'd22628: log10_cal = 16'b0000010101100000;
            15'd22629: log10_cal = 16'b0000010101100000;
            15'd22630: log10_cal = 16'b0000010101100000;
            15'd22631: log10_cal = 16'b0000010101100000;
            15'd22632: log10_cal = 16'b0000010101100000;
            15'd22633: log10_cal = 16'b0000010101100000;
            15'd22634: log10_cal = 16'b0000010101100000;
            15'd22635: log10_cal = 16'b0000010101100000;
            15'd22636: log10_cal = 16'b0000010101100000;
            15'd22637: log10_cal = 16'b0000010101100000;
            15'd22638: log10_cal = 16'b0000010101100000;
            15'd22639: log10_cal = 16'b0000010101100000;
            15'd22640: log10_cal = 16'b0000010101100000;
            15'd22641: log10_cal = 16'b0000010101100000;
            15'd22642: log10_cal = 16'b0000010101100000;
            15'd22643: log10_cal = 16'b0000010101100000;
            15'd22644: log10_cal = 16'b0000010101100000;
            15'd22645: log10_cal = 16'b0000010101100000;
            15'd22646: log10_cal = 16'b0000010101100000;
            15'd22647: log10_cal = 16'b0000010101100000;
            15'd22648: log10_cal = 16'b0000010101100001;
            15'd22649: log10_cal = 16'b0000010101100001;
            15'd22650: log10_cal = 16'b0000010101100001;
            15'd22651: log10_cal = 16'b0000010101100001;
            15'd22652: log10_cal = 16'b0000010101100001;
            15'd22653: log10_cal = 16'b0000010101100001;
            15'd22654: log10_cal = 16'b0000010101100001;
            15'd22655: log10_cal = 16'b0000010101100001;
            15'd22656: log10_cal = 16'b0000010101100001;
            15'd22657: log10_cal = 16'b0000010101100001;
            15'd22658: log10_cal = 16'b0000010101100001;
            15'd22659: log10_cal = 16'b0000010101100001;
            15'd22660: log10_cal = 16'b0000010101100001;
            15'd22661: log10_cal = 16'b0000010101100001;
            15'd22662: log10_cal = 16'b0000010101100001;
            15'd22663: log10_cal = 16'b0000010101100001;
            15'd22664: log10_cal = 16'b0000010101100001;
            15'd22665: log10_cal = 16'b0000010101100001;
            15'd22666: log10_cal = 16'b0000010101100001;
            15'd22667: log10_cal = 16'b0000010101100001;
            15'd22668: log10_cal = 16'b0000010101100001;
            15'd22669: log10_cal = 16'b0000010101100001;
            15'd22670: log10_cal = 16'b0000010101100001;
            15'd22671: log10_cal = 16'b0000010101100001;
            15'd22672: log10_cal = 16'b0000010101100001;
            15'd22673: log10_cal = 16'b0000010101100001;
            15'd22674: log10_cal = 16'b0000010101100001;
            15'd22675: log10_cal = 16'b0000010101100001;
            15'd22676: log10_cal = 16'b0000010101100001;
            15'd22677: log10_cal = 16'b0000010101100001;
            15'd22678: log10_cal = 16'b0000010101100001;
            15'd22679: log10_cal = 16'b0000010101100001;
            15'd22680: log10_cal = 16'b0000010101100001;
            15'd22681: log10_cal = 16'b0000010101100001;
            15'd22682: log10_cal = 16'b0000010101100001;
            15'd22683: log10_cal = 16'b0000010101100001;
            15'd22684: log10_cal = 16'b0000010101100001;
            15'd22685: log10_cal = 16'b0000010101100001;
            15'd22686: log10_cal = 16'b0000010101100001;
            15'd22687: log10_cal = 16'b0000010101100001;
            15'd22688: log10_cal = 16'b0000010101100001;
            15'd22689: log10_cal = 16'b0000010101100001;
            15'd22690: log10_cal = 16'b0000010101100001;
            15'd22691: log10_cal = 16'b0000010101100001;
            15'd22692: log10_cal = 16'b0000010101100001;
            15'd22693: log10_cal = 16'b0000010101100001;
            15'd22694: log10_cal = 16'b0000010101100001;
            15'd22695: log10_cal = 16'b0000010101100001;
            15'd22696: log10_cal = 16'b0000010101100001;
            15'd22697: log10_cal = 16'b0000010101100001;
            15'd22698: log10_cal = 16'b0000010101100001;
            15'd22699: log10_cal = 16'b0000010101100010;
            15'd22700: log10_cal = 16'b0000010101100010;
            15'd22701: log10_cal = 16'b0000010101100010;
            15'd22702: log10_cal = 16'b0000010101100010;
            15'd22703: log10_cal = 16'b0000010101100010;
            15'd22704: log10_cal = 16'b0000010101100010;
            15'd22705: log10_cal = 16'b0000010101100010;
            15'd22706: log10_cal = 16'b0000010101100010;
            15'd22707: log10_cal = 16'b0000010101100010;
            15'd22708: log10_cal = 16'b0000010101100010;
            15'd22709: log10_cal = 16'b0000010101100010;
            15'd22710: log10_cal = 16'b0000010101100010;
            15'd22711: log10_cal = 16'b0000010101100010;
            15'd22712: log10_cal = 16'b0000010101100010;
            15'd22713: log10_cal = 16'b0000010101100010;
            15'd22714: log10_cal = 16'b0000010101100010;
            15'd22715: log10_cal = 16'b0000010101100010;
            15'd22716: log10_cal = 16'b0000010101100010;
            15'd22717: log10_cal = 16'b0000010101100010;
            15'd22718: log10_cal = 16'b0000010101100010;
            15'd22719: log10_cal = 16'b0000010101100010;
            15'd22720: log10_cal = 16'b0000010101100010;
            15'd22721: log10_cal = 16'b0000010101100010;
            15'd22722: log10_cal = 16'b0000010101100010;
            15'd22723: log10_cal = 16'b0000010101100010;
            15'd22724: log10_cal = 16'b0000010101100010;
            15'd22725: log10_cal = 16'b0000010101100010;
            15'd22726: log10_cal = 16'b0000010101100010;
            15'd22727: log10_cal = 16'b0000010101100010;
            15'd22728: log10_cal = 16'b0000010101100010;
            15'd22729: log10_cal = 16'b0000010101100010;
            15'd22730: log10_cal = 16'b0000010101100010;
            15'd22731: log10_cal = 16'b0000010101100010;
            15'd22732: log10_cal = 16'b0000010101100010;
            15'd22733: log10_cal = 16'b0000010101100010;
            15'd22734: log10_cal = 16'b0000010101100010;
            15'd22735: log10_cal = 16'b0000010101100010;
            15'd22736: log10_cal = 16'b0000010101100010;
            15'd22737: log10_cal = 16'b0000010101100010;
            15'd22738: log10_cal = 16'b0000010101100010;
            15'd22739: log10_cal = 16'b0000010101100010;
            15'd22740: log10_cal = 16'b0000010101100010;
            15'd22741: log10_cal = 16'b0000010101100010;
            15'd22742: log10_cal = 16'b0000010101100010;
            15'd22743: log10_cal = 16'b0000010101100010;
            15'd22744: log10_cal = 16'b0000010101100010;
            15'd22745: log10_cal = 16'b0000010101100010;
            15'd22746: log10_cal = 16'b0000010101100010;
            15'd22747: log10_cal = 16'b0000010101100010;
            15'd22748: log10_cal = 16'b0000010101100010;
            15'd22749: log10_cal = 16'b0000010101100010;
            15'd22750: log10_cal = 16'b0000010101100011;
            15'd22751: log10_cal = 16'b0000010101100011;
            15'd22752: log10_cal = 16'b0000010101100011;
            15'd22753: log10_cal = 16'b0000010101100011;
            15'd22754: log10_cal = 16'b0000010101100011;
            15'd22755: log10_cal = 16'b0000010101100011;
            15'd22756: log10_cal = 16'b0000010101100011;
            15'd22757: log10_cal = 16'b0000010101100011;
            15'd22758: log10_cal = 16'b0000010101100011;
            15'd22759: log10_cal = 16'b0000010101100011;
            15'd22760: log10_cal = 16'b0000010101100011;
            15'd22761: log10_cal = 16'b0000010101100011;
            15'd22762: log10_cal = 16'b0000010101100011;
            15'd22763: log10_cal = 16'b0000010101100011;
            15'd22764: log10_cal = 16'b0000010101100011;
            15'd22765: log10_cal = 16'b0000010101100011;
            15'd22766: log10_cal = 16'b0000010101100011;
            15'd22767: log10_cal = 16'b0000010101100011;
            15'd22768: log10_cal = 16'b0000010101100011;
            15'd22769: log10_cal = 16'b0000010101100011;
            15'd22770: log10_cal = 16'b0000010101100011;
            15'd22771: log10_cal = 16'b0000010101100011;
            15'd22772: log10_cal = 16'b0000010101100011;
            15'd22773: log10_cal = 16'b0000010101100011;
            15'd22774: log10_cal = 16'b0000010101100011;
            15'd22775: log10_cal = 16'b0000010101100011;
            15'd22776: log10_cal = 16'b0000010101100011;
            15'd22777: log10_cal = 16'b0000010101100011;
            15'd22778: log10_cal = 16'b0000010101100011;
            15'd22779: log10_cal = 16'b0000010101100011;
            15'd22780: log10_cal = 16'b0000010101100011;
            15'd22781: log10_cal = 16'b0000010101100011;
            15'd22782: log10_cal = 16'b0000010101100011;
            15'd22783: log10_cal = 16'b0000010101100011;
            15'd22784: log10_cal = 16'b0000010101100011;
            15'd22785: log10_cal = 16'b0000010101100011;
            15'd22786: log10_cal = 16'b0000010101100011;
            15'd22787: log10_cal = 16'b0000010101100011;
            15'd22788: log10_cal = 16'b0000010101100011;
            15'd22789: log10_cal = 16'b0000010101100011;
            15'd22790: log10_cal = 16'b0000010101100011;
            15'd22791: log10_cal = 16'b0000010101100011;
            15'd22792: log10_cal = 16'b0000010101100011;
            15'd22793: log10_cal = 16'b0000010101100011;
            15'd22794: log10_cal = 16'b0000010101100011;
            15'd22795: log10_cal = 16'b0000010101100011;
            15'd22796: log10_cal = 16'b0000010101100011;
            15'd22797: log10_cal = 16'b0000010101100011;
            15'd22798: log10_cal = 16'b0000010101100011;
            15'd22799: log10_cal = 16'b0000010101100011;
            15'd22800: log10_cal = 16'b0000010101100011;
            15'd22801: log10_cal = 16'b0000010101100011;
            15'd22802: log10_cal = 16'b0000010101100100;
            15'd22803: log10_cal = 16'b0000010101100100;
            15'd22804: log10_cal = 16'b0000010101100100;
            15'd22805: log10_cal = 16'b0000010101100100;
            15'd22806: log10_cal = 16'b0000010101100100;
            15'd22807: log10_cal = 16'b0000010101100100;
            15'd22808: log10_cal = 16'b0000010101100100;
            15'd22809: log10_cal = 16'b0000010101100100;
            15'd22810: log10_cal = 16'b0000010101100100;
            15'd22811: log10_cal = 16'b0000010101100100;
            15'd22812: log10_cal = 16'b0000010101100100;
            15'd22813: log10_cal = 16'b0000010101100100;
            15'd22814: log10_cal = 16'b0000010101100100;
            15'd22815: log10_cal = 16'b0000010101100100;
            15'd22816: log10_cal = 16'b0000010101100100;
            15'd22817: log10_cal = 16'b0000010101100100;
            15'd22818: log10_cal = 16'b0000010101100100;
            15'd22819: log10_cal = 16'b0000010101100100;
            15'd22820: log10_cal = 16'b0000010101100100;
            15'd22821: log10_cal = 16'b0000010101100100;
            15'd22822: log10_cal = 16'b0000010101100100;
            15'd22823: log10_cal = 16'b0000010101100100;
            15'd22824: log10_cal = 16'b0000010101100100;
            15'd22825: log10_cal = 16'b0000010101100100;
            15'd22826: log10_cal = 16'b0000010101100100;
            15'd22827: log10_cal = 16'b0000010101100100;
            15'd22828: log10_cal = 16'b0000010101100100;
            15'd22829: log10_cal = 16'b0000010101100100;
            15'd22830: log10_cal = 16'b0000010101100100;
            15'd22831: log10_cal = 16'b0000010101100100;
            15'd22832: log10_cal = 16'b0000010101100100;
            15'd22833: log10_cal = 16'b0000010101100100;
            15'd22834: log10_cal = 16'b0000010101100100;
            15'd22835: log10_cal = 16'b0000010101100100;
            15'd22836: log10_cal = 16'b0000010101100100;
            15'd22837: log10_cal = 16'b0000010101100100;
            15'd22838: log10_cal = 16'b0000010101100100;
            15'd22839: log10_cal = 16'b0000010101100100;
            15'd22840: log10_cal = 16'b0000010101100100;
            15'd22841: log10_cal = 16'b0000010101100100;
            15'd22842: log10_cal = 16'b0000010101100100;
            15'd22843: log10_cal = 16'b0000010101100100;
            15'd22844: log10_cal = 16'b0000010101100100;
            15'd22845: log10_cal = 16'b0000010101100100;
            15'd22846: log10_cal = 16'b0000010101100100;
            15'd22847: log10_cal = 16'b0000010101100100;
            15'd22848: log10_cal = 16'b0000010101100100;
            15'd22849: log10_cal = 16'b0000010101100100;
            15'd22850: log10_cal = 16'b0000010101100100;
            15'd22851: log10_cal = 16'b0000010101100100;
            15'd22852: log10_cal = 16'b0000010101100100;
            15'd22853: log10_cal = 16'b0000010101100101;
            15'd22854: log10_cal = 16'b0000010101100101;
            15'd22855: log10_cal = 16'b0000010101100101;
            15'd22856: log10_cal = 16'b0000010101100101;
            15'd22857: log10_cal = 16'b0000010101100101;
            15'd22858: log10_cal = 16'b0000010101100101;
            15'd22859: log10_cal = 16'b0000010101100101;
            15'd22860: log10_cal = 16'b0000010101100101;
            15'd22861: log10_cal = 16'b0000010101100101;
            15'd22862: log10_cal = 16'b0000010101100101;
            15'd22863: log10_cal = 16'b0000010101100101;
            15'd22864: log10_cal = 16'b0000010101100101;
            15'd22865: log10_cal = 16'b0000010101100101;
            15'd22866: log10_cal = 16'b0000010101100101;
            15'd22867: log10_cal = 16'b0000010101100101;
            15'd22868: log10_cal = 16'b0000010101100101;
            15'd22869: log10_cal = 16'b0000010101100101;
            15'd22870: log10_cal = 16'b0000010101100101;
            15'd22871: log10_cal = 16'b0000010101100101;
            15'd22872: log10_cal = 16'b0000010101100101;
            15'd22873: log10_cal = 16'b0000010101100101;
            15'd22874: log10_cal = 16'b0000010101100101;
            15'd22875: log10_cal = 16'b0000010101100101;
            15'd22876: log10_cal = 16'b0000010101100101;
            15'd22877: log10_cal = 16'b0000010101100101;
            15'd22878: log10_cal = 16'b0000010101100101;
            15'd22879: log10_cal = 16'b0000010101100101;
            15'd22880: log10_cal = 16'b0000010101100101;
            15'd22881: log10_cal = 16'b0000010101100101;
            15'd22882: log10_cal = 16'b0000010101100101;
            15'd22883: log10_cal = 16'b0000010101100101;
            15'd22884: log10_cal = 16'b0000010101100101;
            15'd22885: log10_cal = 16'b0000010101100101;
            15'd22886: log10_cal = 16'b0000010101100101;
            15'd22887: log10_cal = 16'b0000010101100101;
            15'd22888: log10_cal = 16'b0000010101100101;
            15'd22889: log10_cal = 16'b0000010101100101;
            15'd22890: log10_cal = 16'b0000010101100101;
            15'd22891: log10_cal = 16'b0000010101100101;
            15'd22892: log10_cal = 16'b0000010101100101;
            15'd22893: log10_cal = 16'b0000010101100101;
            15'd22894: log10_cal = 16'b0000010101100101;
            15'd22895: log10_cal = 16'b0000010101100101;
            15'd22896: log10_cal = 16'b0000010101100101;
            15'd22897: log10_cal = 16'b0000010101100101;
            15'd22898: log10_cal = 16'b0000010101100101;
            15'd22899: log10_cal = 16'b0000010101100101;
            15'd22900: log10_cal = 16'b0000010101100101;
            15'd22901: log10_cal = 16'b0000010101100101;
            15'd22902: log10_cal = 16'b0000010101100101;
            15'd22903: log10_cal = 16'b0000010101100101;
            15'd22904: log10_cal = 16'b0000010101100110;
            15'd22905: log10_cal = 16'b0000010101100110;
            15'd22906: log10_cal = 16'b0000010101100110;
            15'd22907: log10_cal = 16'b0000010101100110;
            15'd22908: log10_cal = 16'b0000010101100110;
            15'd22909: log10_cal = 16'b0000010101100110;
            15'd22910: log10_cal = 16'b0000010101100110;
            15'd22911: log10_cal = 16'b0000010101100110;
            15'd22912: log10_cal = 16'b0000010101100110;
            15'd22913: log10_cal = 16'b0000010101100110;
            15'd22914: log10_cal = 16'b0000010101100110;
            15'd22915: log10_cal = 16'b0000010101100110;
            15'd22916: log10_cal = 16'b0000010101100110;
            15'd22917: log10_cal = 16'b0000010101100110;
            15'd22918: log10_cal = 16'b0000010101100110;
            15'd22919: log10_cal = 16'b0000010101100110;
            15'd22920: log10_cal = 16'b0000010101100110;
            15'd22921: log10_cal = 16'b0000010101100110;
            15'd22922: log10_cal = 16'b0000010101100110;
            15'd22923: log10_cal = 16'b0000010101100110;
            15'd22924: log10_cal = 16'b0000010101100110;
            15'd22925: log10_cal = 16'b0000010101100110;
            15'd22926: log10_cal = 16'b0000010101100110;
            15'd22927: log10_cal = 16'b0000010101100110;
            15'd22928: log10_cal = 16'b0000010101100110;
            15'd22929: log10_cal = 16'b0000010101100110;
            15'd22930: log10_cal = 16'b0000010101100110;
            15'd22931: log10_cal = 16'b0000010101100110;
            15'd22932: log10_cal = 16'b0000010101100110;
            15'd22933: log10_cal = 16'b0000010101100110;
            15'd22934: log10_cal = 16'b0000010101100110;
            15'd22935: log10_cal = 16'b0000010101100110;
            15'd22936: log10_cal = 16'b0000010101100110;
            15'd22937: log10_cal = 16'b0000010101100110;
            15'd22938: log10_cal = 16'b0000010101100110;
            15'd22939: log10_cal = 16'b0000010101100110;
            15'd22940: log10_cal = 16'b0000010101100110;
            15'd22941: log10_cal = 16'b0000010101100110;
            15'd22942: log10_cal = 16'b0000010101100110;
            15'd22943: log10_cal = 16'b0000010101100110;
            15'd22944: log10_cal = 16'b0000010101100110;
            15'd22945: log10_cal = 16'b0000010101100110;
            15'd22946: log10_cal = 16'b0000010101100110;
            15'd22947: log10_cal = 16'b0000010101100110;
            15'd22948: log10_cal = 16'b0000010101100110;
            15'd22949: log10_cal = 16'b0000010101100110;
            15'd22950: log10_cal = 16'b0000010101100110;
            15'd22951: log10_cal = 16'b0000010101100110;
            15'd22952: log10_cal = 16'b0000010101100110;
            15'd22953: log10_cal = 16'b0000010101100110;
            15'd22954: log10_cal = 16'b0000010101100110;
            15'd22955: log10_cal = 16'b0000010101100110;
            15'd22956: log10_cal = 16'b0000010101100111;
            15'd22957: log10_cal = 16'b0000010101100111;
            15'd22958: log10_cal = 16'b0000010101100111;
            15'd22959: log10_cal = 16'b0000010101100111;
            15'd22960: log10_cal = 16'b0000010101100111;
            15'd22961: log10_cal = 16'b0000010101100111;
            15'd22962: log10_cal = 16'b0000010101100111;
            15'd22963: log10_cal = 16'b0000010101100111;
            15'd22964: log10_cal = 16'b0000010101100111;
            15'd22965: log10_cal = 16'b0000010101100111;
            15'd22966: log10_cal = 16'b0000010101100111;
            15'd22967: log10_cal = 16'b0000010101100111;
            15'd22968: log10_cal = 16'b0000010101100111;
            15'd22969: log10_cal = 16'b0000010101100111;
            15'd22970: log10_cal = 16'b0000010101100111;
            15'd22971: log10_cal = 16'b0000010101100111;
            15'd22972: log10_cal = 16'b0000010101100111;
            15'd22973: log10_cal = 16'b0000010101100111;
            15'd22974: log10_cal = 16'b0000010101100111;
            15'd22975: log10_cal = 16'b0000010101100111;
            15'd22976: log10_cal = 16'b0000010101100111;
            15'd22977: log10_cal = 16'b0000010101100111;
            15'd22978: log10_cal = 16'b0000010101100111;
            15'd22979: log10_cal = 16'b0000010101100111;
            15'd22980: log10_cal = 16'b0000010101100111;
            15'd22981: log10_cal = 16'b0000010101100111;
            15'd22982: log10_cal = 16'b0000010101100111;
            15'd22983: log10_cal = 16'b0000010101100111;
            15'd22984: log10_cal = 16'b0000010101100111;
            15'd22985: log10_cal = 16'b0000010101100111;
            15'd22986: log10_cal = 16'b0000010101100111;
            15'd22987: log10_cal = 16'b0000010101100111;
            15'd22988: log10_cal = 16'b0000010101100111;
            15'd22989: log10_cal = 16'b0000010101100111;
            15'd22990: log10_cal = 16'b0000010101100111;
            15'd22991: log10_cal = 16'b0000010101100111;
            15'd22992: log10_cal = 16'b0000010101100111;
            15'd22993: log10_cal = 16'b0000010101100111;
            15'd22994: log10_cal = 16'b0000010101100111;
            15'd22995: log10_cal = 16'b0000010101100111;
            15'd22996: log10_cal = 16'b0000010101100111;
            15'd22997: log10_cal = 16'b0000010101100111;
            15'd22998: log10_cal = 16'b0000010101100111;
            15'd22999: log10_cal = 16'b0000010101100111;
            15'd23000: log10_cal = 16'b0000010101100111;
            15'd23001: log10_cal = 16'b0000010101100111;
            15'd23002: log10_cal = 16'b0000010101100111;
            15'd23003: log10_cal = 16'b0000010101100111;
            15'd23004: log10_cal = 16'b0000010101100111;
            15'd23005: log10_cal = 16'b0000010101100111;
            15'd23006: log10_cal = 16'b0000010101100111;
            15'd23007: log10_cal = 16'b0000010101100111;
            15'd23008: log10_cal = 16'b0000010101101000;
            15'd23009: log10_cal = 16'b0000010101101000;
            15'd23010: log10_cal = 16'b0000010101101000;
            15'd23011: log10_cal = 16'b0000010101101000;
            15'd23012: log10_cal = 16'b0000010101101000;
            15'd23013: log10_cal = 16'b0000010101101000;
            15'd23014: log10_cal = 16'b0000010101101000;
            15'd23015: log10_cal = 16'b0000010101101000;
            15'd23016: log10_cal = 16'b0000010101101000;
            15'd23017: log10_cal = 16'b0000010101101000;
            15'd23018: log10_cal = 16'b0000010101101000;
            15'd23019: log10_cal = 16'b0000010101101000;
            15'd23020: log10_cal = 16'b0000010101101000;
            15'd23021: log10_cal = 16'b0000010101101000;
            15'd23022: log10_cal = 16'b0000010101101000;
            15'd23023: log10_cal = 16'b0000010101101000;
            15'd23024: log10_cal = 16'b0000010101101000;
            15'd23025: log10_cal = 16'b0000010101101000;
            15'd23026: log10_cal = 16'b0000010101101000;
            15'd23027: log10_cal = 16'b0000010101101000;
            15'd23028: log10_cal = 16'b0000010101101000;
            15'd23029: log10_cal = 16'b0000010101101000;
            15'd23030: log10_cal = 16'b0000010101101000;
            15'd23031: log10_cal = 16'b0000010101101000;
            15'd23032: log10_cal = 16'b0000010101101000;
            15'd23033: log10_cal = 16'b0000010101101000;
            15'd23034: log10_cal = 16'b0000010101101000;
            15'd23035: log10_cal = 16'b0000010101101000;
            15'd23036: log10_cal = 16'b0000010101101000;
            15'd23037: log10_cal = 16'b0000010101101000;
            15'd23038: log10_cal = 16'b0000010101101000;
            15'd23039: log10_cal = 16'b0000010101101000;
            15'd23040: log10_cal = 16'b0000010101101000;
            15'd23041: log10_cal = 16'b0000010101101000;
            15'd23042: log10_cal = 16'b0000010101101000;
            15'd23043: log10_cal = 16'b0000010101101000;
            15'd23044: log10_cal = 16'b0000010101101000;
            15'd23045: log10_cal = 16'b0000010101101000;
            15'd23046: log10_cal = 16'b0000010101101000;
            15'd23047: log10_cal = 16'b0000010101101000;
            15'd23048: log10_cal = 16'b0000010101101000;
            15'd23049: log10_cal = 16'b0000010101101000;
            15'd23050: log10_cal = 16'b0000010101101000;
            15'd23051: log10_cal = 16'b0000010101101000;
            15'd23052: log10_cal = 16'b0000010101101000;
            15'd23053: log10_cal = 16'b0000010101101000;
            15'd23054: log10_cal = 16'b0000010101101000;
            15'd23055: log10_cal = 16'b0000010101101000;
            15'd23056: log10_cal = 16'b0000010101101000;
            15'd23057: log10_cal = 16'b0000010101101000;
            15'd23058: log10_cal = 16'b0000010101101000;
            15'd23059: log10_cal = 16'b0000010101101001;
            15'd23060: log10_cal = 16'b0000010101101001;
            15'd23061: log10_cal = 16'b0000010101101001;
            15'd23062: log10_cal = 16'b0000010101101001;
            15'd23063: log10_cal = 16'b0000010101101001;
            15'd23064: log10_cal = 16'b0000010101101001;
            15'd23065: log10_cal = 16'b0000010101101001;
            15'd23066: log10_cal = 16'b0000010101101001;
            15'd23067: log10_cal = 16'b0000010101101001;
            15'd23068: log10_cal = 16'b0000010101101001;
            15'd23069: log10_cal = 16'b0000010101101001;
            15'd23070: log10_cal = 16'b0000010101101001;
            15'd23071: log10_cal = 16'b0000010101101001;
            15'd23072: log10_cal = 16'b0000010101101001;
            15'd23073: log10_cal = 16'b0000010101101001;
            15'd23074: log10_cal = 16'b0000010101101001;
            15'd23075: log10_cal = 16'b0000010101101001;
            15'd23076: log10_cal = 16'b0000010101101001;
            15'd23077: log10_cal = 16'b0000010101101001;
            15'd23078: log10_cal = 16'b0000010101101001;
            15'd23079: log10_cal = 16'b0000010101101001;
            15'd23080: log10_cal = 16'b0000010101101001;
            15'd23081: log10_cal = 16'b0000010101101001;
            15'd23082: log10_cal = 16'b0000010101101001;
            15'd23083: log10_cal = 16'b0000010101101001;
            15'd23084: log10_cal = 16'b0000010101101001;
            15'd23085: log10_cal = 16'b0000010101101001;
            15'd23086: log10_cal = 16'b0000010101101001;
            15'd23087: log10_cal = 16'b0000010101101001;
            15'd23088: log10_cal = 16'b0000010101101001;
            15'd23089: log10_cal = 16'b0000010101101001;
            15'd23090: log10_cal = 16'b0000010101101001;
            15'd23091: log10_cal = 16'b0000010101101001;
            15'd23092: log10_cal = 16'b0000010101101001;
            15'd23093: log10_cal = 16'b0000010101101001;
            15'd23094: log10_cal = 16'b0000010101101001;
            15'd23095: log10_cal = 16'b0000010101101001;
            15'd23096: log10_cal = 16'b0000010101101001;
            15'd23097: log10_cal = 16'b0000010101101001;
            15'd23098: log10_cal = 16'b0000010101101001;
            15'd23099: log10_cal = 16'b0000010101101001;
            15'd23100: log10_cal = 16'b0000010101101001;
            15'd23101: log10_cal = 16'b0000010101101001;
            15'd23102: log10_cal = 16'b0000010101101001;
            15'd23103: log10_cal = 16'b0000010101101001;
            15'd23104: log10_cal = 16'b0000010101101001;
            15'd23105: log10_cal = 16'b0000010101101001;
            15'd23106: log10_cal = 16'b0000010101101001;
            15'd23107: log10_cal = 16'b0000010101101001;
            15'd23108: log10_cal = 16'b0000010101101001;
            15'd23109: log10_cal = 16'b0000010101101001;
            15'd23110: log10_cal = 16'b0000010101101001;
            15'd23111: log10_cal = 16'b0000010101101010;
            15'd23112: log10_cal = 16'b0000010101101010;
            15'd23113: log10_cal = 16'b0000010101101010;
            15'd23114: log10_cal = 16'b0000010101101010;
            15'd23115: log10_cal = 16'b0000010101101010;
            15'd23116: log10_cal = 16'b0000010101101010;
            15'd23117: log10_cal = 16'b0000010101101010;
            15'd23118: log10_cal = 16'b0000010101101010;
            15'd23119: log10_cal = 16'b0000010101101010;
            15'd23120: log10_cal = 16'b0000010101101010;
            15'd23121: log10_cal = 16'b0000010101101010;
            15'd23122: log10_cal = 16'b0000010101101010;
            15'd23123: log10_cal = 16'b0000010101101010;
            15'd23124: log10_cal = 16'b0000010101101010;
            15'd23125: log10_cal = 16'b0000010101101010;
            15'd23126: log10_cal = 16'b0000010101101010;
            15'd23127: log10_cal = 16'b0000010101101010;
            15'd23128: log10_cal = 16'b0000010101101010;
            15'd23129: log10_cal = 16'b0000010101101010;
            15'd23130: log10_cal = 16'b0000010101101010;
            15'd23131: log10_cal = 16'b0000010101101010;
            15'd23132: log10_cal = 16'b0000010101101010;
            15'd23133: log10_cal = 16'b0000010101101010;
            15'd23134: log10_cal = 16'b0000010101101010;
            15'd23135: log10_cal = 16'b0000010101101010;
            15'd23136: log10_cal = 16'b0000010101101010;
            15'd23137: log10_cal = 16'b0000010101101010;
            15'd23138: log10_cal = 16'b0000010101101010;
            15'd23139: log10_cal = 16'b0000010101101010;
            15'd23140: log10_cal = 16'b0000010101101010;
            15'd23141: log10_cal = 16'b0000010101101010;
            15'd23142: log10_cal = 16'b0000010101101010;
            15'd23143: log10_cal = 16'b0000010101101010;
            15'd23144: log10_cal = 16'b0000010101101010;
            15'd23145: log10_cal = 16'b0000010101101010;
            15'd23146: log10_cal = 16'b0000010101101010;
            15'd23147: log10_cal = 16'b0000010101101010;
            15'd23148: log10_cal = 16'b0000010101101010;
            15'd23149: log10_cal = 16'b0000010101101010;
            15'd23150: log10_cal = 16'b0000010101101010;
            15'd23151: log10_cal = 16'b0000010101101010;
            15'd23152: log10_cal = 16'b0000010101101010;
            15'd23153: log10_cal = 16'b0000010101101010;
            15'd23154: log10_cal = 16'b0000010101101010;
            15'd23155: log10_cal = 16'b0000010101101010;
            15'd23156: log10_cal = 16'b0000010101101010;
            15'd23157: log10_cal = 16'b0000010101101010;
            15'd23158: log10_cal = 16'b0000010101101010;
            15'd23159: log10_cal = 16'b0000010101101010;
            15'd23160: log10_cal = 16'b0000010101101010;
            15'd23161: log10_cal = 16'b0000010101101010;
            15'd23162: log10_cal = 16'b0000010101101010;
            15'd23163: log10_cal = 16'b0000010101101011;
            15'd23164: log10_cal = 16'b0000010101101011;
            15'd23165: log10_cal = 16'b0000010101101011;
            15'd23166: log10_cal = 16'b0000010101101011;
            15'd23167: log10_cal = 16'b0000010101101011;
            15'd23168: log10_cal = 16'b0000010101101011;
            15'd23169: log10_cal = 16'b0000010101101011;
            15'd23170: log10_cal = 16'b0000010101101011;
            15'd23171: log10_cal = 16'b0000010101101011;
            15'd23172: log10_cal = 16'b0000010101101011;
            15'd23173: log10_cal = 16'b0000010101101011;
            15'd23174: log10_cal = 16'b0000010101101011;
            15'd23175: log10_cal = 16'b0000010101101011;
            15'd23176: log10_cal = 16'b0000010101101011;
            15'd23177: log10_cal = 16'b0000010101101011;
            15'd23178: log10_cal = 16'b0000010101101011;
            15'd23179: log10_cal = 16'b0000010101101011;
            15'd23180: log10_cal = 16'b0000010101101011;
            15'd23181: log10_cal = 16'b0000010101101011;
            15'd23182: log10_cal = 16'b0000010101101011;
            15'd23183: log10_cal = 16'b0000010101101011;
            15'd23184: log10_cal = 16'b0000010101101011;
            15'd23185: log10_cal = 16'b0000010101101011;
            15'd23186: log10_cal = 16'b0000010101101011;
            15'd23187: log10_cal = 16'b0000010101101011;
            15'd23188: log10_cal = 16'b0000010101101011;
            15'd23189: log10_cal = 16'b0000010101101011;
            15'd23190: log10_cal = 16'b0000010101101011;
            15'd23191: log10_cal = 16'b0000010101101011;
            15'd23192: log10_cal = 16'b0000010101101011;
            15'd23193: log10_cal = 16'b0000010101101011;
            15'd23194: log10_cal = 16'b0000010101101011;
            15'd23195: log10_cal = 16'b0000010101101011;
            15'd23196: log10_cal = 16'b0000010101101011;
            15'd23197: log10_cal = 16'b0000010101101011;
            15'd23198: log10_cal = 16'b0000010101101011;
            15'd23199: log10_cal = 16'b0000010101101011;
            15'd23200: log10_cal = 16'b0000010101101011;
            15'd23201: log10_cal = 16'b0000010101101011;
            15'd23202: log10_cal = 16'b0000010101101011;
            15'd23203: log10_cal = 16'b0000010101101011;
            15'd23204: log10_cal = 16'b0000010101101011;
            15'd23205: log10_cal = 16'b0000010101101011;
            15'd23206: log10_cal = 16'b0000010101101011;
            15'd23207: log10_cal = 16'b0000010101101011;
            15'd23208: log10_cal = 16'b0000010101101011;
            15'd23209: log10_cal = 16'b0000010101101011;
            15'd23210: log10_cal = 16'b0000010101101011;
            15'd23211: log10_cal = 16'b0000010101101011;
            15'd23212: log10_cal = 16'b0000010101101011;
            15'd23213: log10_cal = 16'b0000010101101011;
            15'd23214: log10_cal = 16'b0000010101101011;
            15'd23215: log10_cal = 16'b0000010101101011;
            15'd23216: log10_cal = 16'b0000010101101100;
            15'd23217: log10_cal = 16'b0000010101101100;
            15'd23218: log10_cal = 16'b0000010101101100;
            15'd23219: log10_cal = 16'b0000010101101100;
            15'd23220: log10_cal = 16'b0000010101101100;
            15'd23221: log10_cal = 16'b0000010101101100;
            15'd23222: log10_cal = 16'b0000010101101100;
            15'd23223: log10_cal = 16'b0000010101101100;
            15'd23224: log10_cal = 16'b0000010101101100;
            15'd23225: log10_cal = 16'b0000010101101100;
            15'd23226: log10_cal = 16'b0000010101101100;
            15'd23227: log10_cal = 16'b0000010101101100;
            15'd23228: log10_cal = 16'b0000010101101100;
            15'd23229: log10_cal = 16'b0000010101101100;
            15'd23230: log10_cal = 16'b0000010101101100;
            15'd23231: log10_cal = 16'b0000010101101100;
            15'd23232: log10_cal = 16'b0000010101101100;
            15'd23233: log10_cal = 16'b0000010101101100;
            15'd23234: log10_cal = 16'b0000010101101100;
            15'd23235: log10_cal = 16'b0000010101101100;
            15'd23236: log10_cal = 16'b0000010101101100;
            15'd23237: log10_cal = 16'b0000010101101100;
            15'd23238: log10_cal = 16'b0000010101101100;
            15'd23239: log10_cal = 16'b0000010101101100;
            15'd23240: log10_cal = 16'b0000010101101100;
            15'd23241: log10_cal = 16'b0000010101101100;
            15'd23242: log10_cal = 16'b0000010101101100;
            15'd23243: log10_cal = 16'b0000010101101100;
            15'd23244: log10_cal = 16'b0000010101101100;
            15'd23245: log10_cal = 16'b0000010101101100;
            15'd23246: log10_cal = 16'b0000010101101100;
            15'd23247: log10_cal = 16'b0000010101101100;
            15'd23248: log10_cal = 16'b0000010101101100;
            15'd23249: log10_cal = 16'b0000010101101100;
            15'd23250: log10_cal = 16'b0000010101101100;
            15'd23251: log10_cal = 16'b0000010101101100;
            15'd23252: log10_cal = 16'b0000010101101100;
            15'd23253: log10_cal = 16'b0000010101101100;
            15'd23254: log10_cal = 16'b0000010101101100;
            15'd23255: log10_cal = 16'b0000010101101100;
            15'd23256: log10_cal = 16'b0000010101101100;
            15'd23257: log10_cal = 16'b0000010101101100;
            15'd23258: log10_cal = 16'b0000010101101100;
            15'd23259: log10_cal = 16'b0000010101101100;
            15'd23260: log10_cal = 16'b0000010101101100;
            15'd23261: log10_cal = 16'b0000010101101100;
            15'd23262: log10_cal = 16'b0000010101101100;
            15'd23263: log10_cal = 16'b0000010101101100;
            15'd23264: log10_cal = 16'b0000010101101100;
            15'd23265: log10_cal = 16'b0000010101101100;
            15'd23266: log10_cal = 16'b0000010101101100;
            15'd23267: log10_cal = 16'b0000010101101100;
            15'd23268: log10_cal = 16'b0000010101101101;
            15'd23269: log10_cal = 16'b0000010101101101;
            15'd23270: log10_cal = 16'b0000010101101101;
            15'd23271: log10_cal = 16'b0000010101101101;
            15'd23272: log10_cal = 16'b0000010101101101;
            15'd23273: log10_cal = 16'b0000010101101101;
            15'd23274: log10_cal = 16'b0000010101101101;
            15'd23275: log10_cal = 16'b0000010101101101;
            15'd23276: log10_cal = 16'b0000010101101101;
            15'd23277: log10_cal = 16'b0000010101101101;
            15'd23278: log10_cal = 16'b0000010101101101;
            15'd23279: log10_cal = 16'b0000010101101101;
            15'd23280: log10_cal = 16'b0000010101101101;
            15'd23281: log10_cal = 16'b0000010101101101;
            15'd23282: log10_cal = 16'b0000010101101101;
            15'd23283: log10_cal = 16'b0000010101101101;
            15'd23284: log10_cal = 16'b0000010101101101;
            15'd23285: log10_cal = 16'b0000010101101101;
            15'd23286: log10_cal = 16'b0000010101101101;
            15'd23287: log10_cal = 16'b0000010101101101;
            15'd23288: log10_cal = 16'b0000010101101101;
            15'd23289: log10_cal = 16'b0000010101101101;
            15'd23290: log10_cal = 16'b0000010101101101;
            15'd23291: log10_cal = 16'b0000010101101101;
            15'd23292: log10_cal = 16'b0000010101101101;
            15'd23293: log10_cal = 16'b0000010101101101;
            15'd23294: log10_cal = 16'b0000010101101101;
            15'd23295: log10_cal = 16'b0000010101101101;
            15'd23296: log10_cal = 16'b0000010101101101;
            15'd23297: log10_cal = 16'b0000010101101101;
            15'd23298: log10_cal = 16'b0000010101101101;
            15'd23299: log10_cal = 16'b0000010101101101;
            15'd23300: log10_cal = 16'b0000010101101101;
            15'd23301: log10_cal = 16'b0000010101101101;
            15'd23302: log10_cal = 16'b0000010101101101;
            15'd23303: log10_cal = 16'b0000010101101101;
            15'd23304: log10_cal = 16'b0000010101101101;
            15'd23305: log10_cal = 16'b0000010101101101;
            15'd23306: log10_cal = 16'b0000010101101101;
            15'd23307: log10_cal = 16'b0000010101101101;
            15'd23308: log10_cal = 16'b0000010101101101;
            15'd23309: log10_cal = 16'b0000010101101101;
            15'd23310: log10_cal = 16'b0000010101101101;
            15'd23311: log10_cal = 16'b0000010101101101;
            15'd23312: log10_cal = 16'b0000010101101101;
            15'd23313: log10_cal = 16'b0000010101101101;
            15'd23314: log10_cal = 16'b0000010101101101;
            15'd23315: log10_cal = 16'b0000010101101101;
            15'd23316: log10_cal = 16'b0000010101101101;
            15'd23317: log10_cal = 16'b0000010101101101;
            15'd23318: log10_cal = 16'b0000010101101101;
            15'd23319: log10_cal = 16'b0000010101101101;
            15'd23320: log10_cal = 16'b0000010101101110;
            15'd23321: log10_cal = 16'b0000010101101110;
            15'd23322: log10_cal = 16'b0000010101101110;
            15'd23323: log10_cal = 16'b0000010101101110;
            15'd23324: log10_cal = 16'b0000010101101110;
            15'd23325: log10_cal = 16'b0000010101101110;
            15'd23326: log10_cal = 16'b0000010101101110;
            15'd23327: log10_cal = 16'b0000010101101110;
            15'd23328: log10_cal = 16'b0000010101101110;
            15'd23329: log10_cal = 16'b0000010101101110;
            15'd23330: log10_cal = 16'b0000010101101110;
            15'd23331: log10_cal = 16'b0000010101101110;
            15'd23332: log10_cal = 16'b0000010101101110;
            15'd23333: log10_cal = 16'b0000010101101110;
            15'd23334: log10_cal = 16'b0000010101101110;
            15'd23335: log10_cal = 16'b0000010101101110;
            15'd23336: log10_cal = 16'b0000010101101110;
            15'd23337: log10_cal = 16'b0000010101101110;
            15'd23338: log10_cal = 16'b0000010101101110;
            15'd23339: log10_cal = 16'b0000010101101110;
            15'd23340: log10_cal = 16'b0000010101101110;
            15'd23341: log10_cal = 16'b0000010101101110;
            15'd23342: log10_cal = 16'b0000010101101110;
            15'd23343: log10_cal = 16'b0000010101101110;
            15'd23344: log10_cal = 16'b0000010101101110;
            15'd23345: log10_cal = 16'b0000010101101110;
            15'd23346: log10_cal = 16'b0000010101101110;
            15'd23347: log10_cal = 16'b0000010101101110;
            15'd23348: log10_cal = 16'b0000010101101110;
            15'd23349: log10_cal = 16'b0000010101101110;
            15'd23350: log10_cal = 16'b0000010101101110;
            15'd23351: log10_cal = 16'b0000010101101110;
            15'd23352: log10_cal = 16'b0000010101101110;
            15'd23353: log10_cal = 16'b0000010101101110;
            15'd23354: log10_cal = 16'b0000010101101110;
            15'd23355: log10_cal = 16'b0000010101101110;
            15'd23356: log10_cal = 16'b0000010101101110;
            15'd23357: log10_cal = 16'b0000010101101110;
            15'd23358: log10_cal = 16'b0000010101101110;
            15'd23359: log10_cal = 16'b0000010101101110;
            15'd23360: log10_cal = 16'b0000010101101110;
            15'd23361: log10_cal = 16'b0000010101101110;
            15'd23362: log10_cal = 16'b0000010101101110;
            15'd23363: log10_cal = 16'b0000010101101110;
            15'd23364: log10_cal = 16'b0000010101101110;
            15'd23365: log10_cal = 16'b0000010101101110;
            15'd23366: log10_cal = 16'b0000010101101110;
            15'd23367: log10_cal = 16'b0000010101101110;
            15'd23368: log10_cal = 16'b0000010101101110;
            15'd23369: log10_cal = 16'b0000010101101110;
            15'd23370: log10_cal = 16'b0000010101101110;
            15'd23371: log10_cal = 16'b0000010101101110;
            15'd23372: log10_cal = 16'b0000010101101110;
            15'd23373: log10_cal = 16'b0000010101101111;
            15'd23374: log10_cal = 16'b0000010101101111;
            15'd23375: log10_cal = 16'b0000010101101111;
            15'd23376: log10_cal = 16'b0000010101101111;
            15'd23377: log10_cal = 16'b0000010101101111;
            15'd23378: log10_cal = 16'b0000010101101111;
            15'd23379: log10_cal = 16'b0000010101101111;
            15'd23380: log10_cal = 16'b0000010101101111;
            15'd23381: log10_cal = 16'b0000010101101111;
            15'd23382: log10_cal = 16'b0000010101101111;
            15'd23383: log10_cal = 16'b0000010101101111;
            15'd23384: log10_cal = 16'b0000010101101111;
            15'd23385: log10_cal = 16'b0000010101101111;
            15'd23386: log10_cal = 16'b0000010101101111;
            15'd23387: log10_cal = 16'b0000010101101111;
            15'd23388: log10_cal = 16'b0000010101101111;
            15'd23389: log10_cal = 16'b0000010101101111;
            15'd23390: log10_cal = 16'b0000010101101111;
            15'd23391: log10_cal = 16'b0000010101101111;
            15'd23392: log10_cal = 16'b0000010101101111;
            15'd23393: log10_cal = 16'b0000010101101111;
            15'd23394: log10_cal = 16'b0000010101101111;
            15'd23395: log10_cal = 16'b0000010101101111;
            15'd23396: log10_cal = 16'b0000010101101111;
            15'd23397: log10_cal = 16'b0000010101101111;
            15'd23398: log10_cal = 16'b0000010101101111;
            15'd23399: log10_cal = 16'b0000010101101111;
            15'd23400: log10_cal = 16'b0000010101101111;
            15'd23401: log10_cal = 16'b0000010101101111;
            15'd23402: log10_cal = 16'b0000010101101111;
            15'd23403: log10_cal = 16'b0000010101101111;
            15'd23404: log10_cal = 16'b0000010101101111;
            15'd23405: log10_cal = 16'b0000010101101111;
            15'd23406: log10_cal = 16'b0000010101101111;
            15'd23407: log10_cal = 16'b0000010101101111;
            15'd23408: log10_cal = 16'b0000010101101111;
            15'd23409: log10_cal = 16'b0000010101101111;
            15'd23410: log10_cal = 16'b0000010101101111;
            15'd23411: log10_cal = 16'b0000010101101111;
            15'd23412: log10_cal = 16'b0000010101101111;
            15'd23413: log10_cal = 16'b0000010101101111;
            15'd23414: log10_cal = 16'b0000010101101111;
            15'd23415: log10_cal = 16'b0000010101101111;
            15'd23416: log10_cal = 16'b0000010101101111;
            15'd23417: log10_cal = 16'b0000010101101111;
            15'd23418: log10_cal = 16'b0000010101101111;
            15'd23419: log10_cal = 16'b0000010101101111;
            15'd23420: log10_cal = 16'b0000010101101111;
            15'd23421: log10_cal = 16'b0000010101101111;
            15'd23422: log10_cal = 16'b0000010101101111;
            15'd23423: log10_cal = 16'b0000010101101111;
            15'd23424: log10_cal = 16'b0000010101101111;
            15'd23425: log10_cal = 16'b0000010101110000;
            15'd23426: log10_cal = 16'b0000010101110000;
            15'd23427: log10_cal = 16'b0000010101110000;
            15'd23428: log10_cal = 16'b0000010101110000;
            15'd23429: log10_cal = 16'b0000010101110000;
            15'd23430: log10_cal = 16'b0000010101110000;
            15'd23431: log10_cal = 16'b0000010101110000;
            15'd23432: log10_cal = 16'b0000010101110000;
            15'd23433: log10_cal = 16'b0000010101110000;
            15'd23434: log10_cal = 16'b0000010101110000;
            15'd23435: log10_cal = 16'b0000010101110000;
            15'd23436: log10_cal = 16'b0000010101110000;
            15'd23437: log10_cal = 16'b0000010101110000;
            15'd23438: log10_cal = 16'b0000010101110000;
            15'd23439: log10_cal = 16'b0000010101110000;
            15'd23440: log10_cal = 16'b0000010101110000;
            15'd23441: log10_cal = 16'b0000010101110000;
            15'd23442: log10_cal = 16'b0000010101110000;
            15'd23443: log10_cal = 16'b0000010101110000;
            15'd23444: log10_cal = 16'b0000010101110000;
            15'd23445: log10_cal = 16'b0000010101110000;
            15'd23446: log10_cal = 16'b0000010101110000;
            15'd23447: log10_cal = 16'b0000010101110000;
            15'd23448: log10_cal = 16'b0000010101110000;
            15'd23449: log10_cal = 16'b0000010101110000;
            15'd23450: log10_cal = 16'b0000010101110000;
            15'd23451: log10_cal = 16'b0000010101110000;
            15'd23452: log10_cal = 16'b0000010101110000;
            15'd23453: log10_cal = 16'b0000010101110000;
            15'd23454: log10_cal = 16'b0000010101110000;
            15'd23455: log10_cal = 16'b0000010101110000;
            15'd23456: log10_cal = 16'b0000010101110000;
            15'd23457: log10_cal = 16'b0000010101110000;
            15'd23458: log10_cal = 16'b0000010101110000;
            15'd23459: log10_cal = 16'b0000010101110000;
            15'd23460: log10_cal = 16'b0000010101110000;
            15'd23461: log10_cal = 16'b0000010101110000;
            15'd23462: log10_cal = 16'b0000010101110000;
            15'd23463: log10_cal = 16'b0000010101110000;
            15'd23464: log10_cal = 16'b0000010101110000;
            15'd23465: log10_cal = 16'b0000010101110000;
            15'd23466: log10_cal = 16'b0000010101110000;
            15'd23467: log10_cal = 16'b0000010101110000;
            15'd23468: log10_cal = 16'b0000010101110000;
            15'd23469: log10_cal = 16'b0000010101110000;
            15'd23470: log10_cal = 16'b0000010101110000;
            15'd23471: log10_cal = 16'b0000010101110000;
            15'd23472: log10_cal = 16'b0000010101110000;
            15'd23473: log10_cal = 16'b0000010101110000;
            15'd23474: log10_cal = 16'b0000010101110000;
            15'd23475: log10_cal = 16'b0000010101110000;
            15'd23476: log10_cal = 16'b0000010101110000;
            15'd23477: log10_cal = 16'b0000010101110000;
            15'd23478: log10_cal = 16'b0000010101110001;
            15'd23479: log10_cal = 16'b0000010101110001;
            15'd23480: log10_cal = 16'b0000010101110001;
            15'd23481: log10_cal = 16'b0000010101110001;
            15'd23482: log10_cal = 16'b0000010101110001;
            15'd23483: log10_cal = 16'b0000010101110001;
            15'd23484: log10_cal = 16'b0000010101110001;
            15'd23485: log10_cal = 16'b0000010101110001;
            15'd23486: log10_cal = 16'b0000010101110001;
            15'd23487: log10_cal = 16'b0000010101110001;
            15'd23488: log10_cal = 16'b0000010101110001;
            15'd23489: log10_cal = 16'b0000010101110001;
            15'd23490: log10_cal = 16'b0000010101110001;
            15'd23491: log10_cal = 16'b0000010101110001;
            15'd23492: log10_cal = 16'b0000010101110001;
            15'd23493: log10_cal = 16'b0000010101110001;
            15'd23494: log10_cal = 16'b0000010101110001;
            15'd23495: log10_cal = 16'b0000010101110001;
            15'd23496: log10_cal = 16'b0000010101110001;
            15'd23497: log10_cal = 16'b0000010101110001;
            15'd23498: log10_cal = 16'b0000010101110001;
            15'd23499: log10_cal = 16'b0000010101110001;
            15'd23500: log10_cal = 16'b0000010101110001;
            15'd23501: log10_cal = 16'b0000010101110001;
            15'd23502: log10_cal = 16'b0000010101110001;
            15'd23503: log10_cal = 16'b0000010101110001;
            15'd23504: log10_cal = 16'b0000010101110001;
            15'd23505: log10_cal = 16'b0000010101110001;
            15'd23506: log10_cal = 16'b0000010101110001;
            15'd23507: log10_cal = 16'b0000010101110001;
            15'd23508: log10_cal = 16'b0000010101110001;
            15'd23509: log10_cal = 16'b0000010101110001;
            15'd23510: log10_cal = 16'b0000010101110001;
            15'd23511: log10_cal = 16'b0000010101110001;
            15'd23512: log10_cal = 16'b0000010101110001;
            15'd23513: log10_cal = 16'b0000010101110001;
            15'd23514: log10_cal = 16'b0000010101110001;
            15'd23515: log10_cal = 16'b0000010101110001;
            15'd23516: log10_cal = 16'b0000010101110001;
            15'd23517: log10_cal = 16'b0000010101110001;
            15'd23518: log10_cal = 16'b0000010101110001;
            15'd23519: log10_cal = 16'b0000010101110001;
            15'd23520: log10_cal = 16'b0000010101110001;
            15'd23521: log10_cal = 16'b0000010101110001;
            15'd23522: log10_cal = 16'b0000010101110001;
            15'd23523: log10_cal = 16'b0000010101110001;
            15'd23524: log10_cal = 16'b0000010101110001;
            15'd23525: log10_cal = 16'b0000010101110001;
            15'd23526: log10_cal = 16'b0000010101110001;
            15'd23527: log10_cal = 16'b0000010101110001;
            15'd23528: log10_cal = 16'b0000010101110001;
            15'd23529: log10_cal = 16'b0000010101110001;
            15'd23530: log10_cal = 16'b0000010101110001;
            15'd23531: log10_cal = 16'b0000010101110010;
            15'd23532: log10_cal = 16'b0000010101110010;
            15'd23533: log10_cal = 16'b0000010101110010;
            15'd23534: log10_cal = 16'b0000010101110010;
            15'd23535: log10_cal = 16'b0000010101110010;
            15'd23536: log10_cal = 16'b0000010101110010;
            15'd23537: log10_cal = 16'b0000010101110010;
            15'd23538: log10_cal = 16'b0000010101110010;
            15'd23539: log10_cal = 16'b0000010101110010;
            15'd23540: log10_cal = 16'b0000010101110010;
            15'd23541: log10_cal = 16'b0000010101110010;
            15'd23542: log10_cal = 16'b0000010101110010;
            15'd23543: log10_cal = 16'b0000010101110010;
            15'd23544: log10_cal = 16'b0000010101110010;
            15'd23545: log10_cal = 16'b0000010101110010;
            15'd23546: log10_cal = 16'b0000010101110010;
            15'd23547: log10_cal = 16'b0000010101110010;
            15'd23548: log10_cal = 16'b0000010101110010;
            15'd23549: log10_cal = 16'b0000010101110010;
            15'd23550: log10_cal = 16'b0000010101110010;
            15'd23551: log10_cal = 16'b0000010101110010;
            15'd23552: log10_cal = 16'b0000010101110010;
            15'd23553: log10_cal = 16'b0000010101110010;
            15'd23554: log10_cal = 16'b0000010101110010;
            15'd23555: log10_cal = 16'b0000010101110010;
            15'd23556: log10_cal = 16'b0000010101110010;
            15'd23557: log10_cal = 16'b0000010101110010;
            15'd23558: log10_cal = 16'b0000010101110010;
            15'd23559: log10_cal = 16'b0000010101110010;
            15'd23560: log10_cal = 16'b0000010101110010;
            15'd23561: log10_cal = 16'b0000010101110010;
            15'd23562: log10_cal = 16'b0000010101110010;
            15'd23563: log10_cal = 16'b0000010101110010;
            15'd23564: log10_cal = 16'b0000010101110010;
            15'd23565: log10_cal = 16'b0000010101110010;
            15'd23566: log10_cal = 16'b0000010101110010;
            15'd23567: log10_cal = 16'b0000010101110010;
            15'd23568: log10_cal = 16'b0000010101110010;
            15'd23569: log10_cal = 16'b0000010101110010;
            15'd23570: log10_cal = 16'b0000010101110010;
            15'd23571: log10_cal = 16'b0000010101110010;
            15'd23572: log10_cal = 16'b0000010101110010;
            15'd23573: log10_cal = 16'b0000010101110010;
            15'd23574: log10_cal = 16'b0000010101110010;
            15'd23575: log10_cal = 16'b0000010101110010;
            15'd23576: log10_cal = 16'b0000010101110010;
            15'd23577: log10_cal = 16'b0000010101110010;
            15'd23578: log10_cal = 16'b0000010101110010;
            15'd23579: log10_cal = 16'b0000010101110010;
            15'd23580: log10_cal = 16'b0000010101110010;
            15'd23581: log10_cal = 16'b0000010101110010;
            15'd23582: log10_cal = 16'b0000010101110010;
            15'd23583: log10_cal = 16'b0000010101110010;
            15'd23584: log10_cal = 16'b0000010101110011;
            15'd23585: log10_cal = 16'b0000010101110011;
            15'd23586: log10_cal = 16'b0000010101110011;
            15'd23587: log10_cal = 16'b0000010101110011;
            15'd23588: log10_cal = 16'b0000010101110011;
            15'd23589: log10_cal = 16'b0000010101110011;
            15'd23590: log10_cal = 16'b0000010101110011;
            15'd23591: log10_cal = 16'b0000010101110011;
            15'd23592: log10_cal = 16'b0000010101110011;
            15'd23593: log10_cal = 16'b0000010101110011;
            15'd23594: log10_cal = 16'b0000010101110011;
            15'd23595: log10_cal = 16'b0000010101110011;
            15'd23596: log10_cal = 16'b0000010101110011;
            15'd23597: log10_cal = 16'b0000010101110011;
            15'd23598: log10_cal = 16'b0000010101110011;
            15'd23599: log10_cal = 16'b0000010101110011;
            15'd23600: log10_cal = 16'b0000010101110011;
            15'd23601: log10_cal = 16'b0000010101110011;
            15'd23602: log10_cal = 16'b0000010101110011;
            15'd23603: log10_cal = 16'b0000010101110011;
            15'd23604: log10_cal = 16'b0000010101110011;
            15'd23605: log10_cal = 16'b0000010101110011;
            15'd23606: log10_cal = 16'b0000010101110011;
            15'd23607: log10_cal = 16'b0000010101110011;
            15'd23608: log10_cal = 16'b0000010101110011;
            15'd23609: log10_cal = 16'b0000010101110011;
            15'd23610: log10_cal = 16'b0000010101110011;
            15'd23611: log10_cal = 16'b0000010101110011;
            15'd23612: log10_cal = 16'b0000010101110011;
            15'd23613: log10_cal = 16'b0000010101110011;
            15'd23614: log10_cal = 16'b0000010101110011;
            15'd23615: log10_cal = 16'b0000010101110011;
            15'd23616: log10_cal = 16'b0000010101110011;
            15'd23617: log10_cal = 16'b0000010101110011;
            15'd23618: log10_cal = 16'b0000010101110011;
            15'd23619: log10_cal = 16'b0000010101110011;
            15'd23620: log10_cal = 16'b0000010101110011;
            15'd23621: log10_cal = 16'b0000010101110011;
            15'd23622: log10_cal = 16'b0000010101110011;
            15'd23623: log10_cal = 16'b0000010101110011;
            15'd23624: log10_cal = 16'b0000010101110011;
            15'd23625: log10_cal = 16'b0000010101110011;
            15'd23626: log10_cal = 16'b0000010101110011;
            15'd23627: log10_cal = 16'b0000010101110011;
            15'd23628: log10_cal = 16'b0000010101110011;
            15'd23629: log10_cal = 16'b0000010101110011;
            15'd23630: log10_cal = 16'b0000010101110011;
            15'd23631: log10_cal = 16'b0000010101110011;
            15'd23632: log10_cal = 16'b0000010101110011;
            15'd23633: log10_cal = 16'b0000010101110011;
            15'd23634: log10_cal = 16'b0000010101110011;
            15'd23635: log10_cal = 16'b0000010101110011;
            15'd23636: log10_cal = 16'b0000010101110011;
            15'd23637: log10_cal = 16'b0000010101110100;
            15'd23638: log10_cal = 16'b0000010101110100;
            15'd23639: log10_cal = 16'b0000010101110100;
            15'd23640: log10_cal = 16'b0000010101110100;
            15'd23641: log10_cal = 16'b0000010101110100;
            15'd23642: log10_cal = 16'b0000010101110100;
            15'd23643: log10_cal = 16'b0000010101110100;
            15'd23644: log10_cal = 16'b0000010101110100;
            15'd23645: log10_cal = 16'b0000010101110100;
            15'd23646: log10_cal = 16'b0000010101110100;
            15'd23647: log10_cal = 16'b0000010101110100;
            15'd23648: log10_cal = 16'b0000010101110100;
            15'd23649: log10_cal = 16'b0000010101110100;
            15'd23650: log10_cal = 16'b0000010101110100;
            15'd23651: log10_cal = 16'b0000010101110100;
            15'd23652: log10_cal = 16'b0000010101110100;
            15'd23653: log10_cal = 16'b0000010101110100;
            15'd23654: log10_cal = 16'b0000010101110100;
            15'd23655: log10_cal = 16'b0000010101110100;
            15'd23656: log10_cal = 16'b0000010101110100;
            15'd23657: log10_cal = 16'b0000010101110100;
            15'd23658: log10_cal = 16'b0000010101110100;
            15'd23659: log10_cal = 16'b0000010101110100;
            15'd23660: log10_cal = 16'b0000010101110100;
            15'd23661: log10_cal = 16'b0000010101110100;
            15'd23662: log10_cal = 16'b0000010101110100;
            15'd23663: log10_cal = 16'b0000010101110100;
            15'd23664: log10_cal = 16'b0000010101110100;
            15'd23665: log10_cal = 16'b0000010101110100;
            15'd23666: log10_cal = 16'b0000010101110100;
            15'd23667: log10_cal = 16'b0000010101110100;
            15'd23668: log10_cal = 16'b0000010101110100;
            15'd23669: log10_cal = 16'b0000010101110100;
            15'd23670: log10_cal = 16'b0000010101110100;
            15'd23671: log10_cal = 16'b0000010101110100;
            15'd23672: log10_cal = 16'b0000010101110100;
            15'd23673: log10_cal = 16'b0000010101110100;
            15'd23674: log10_cal = 16'b0000010101110100;
            15'd23675: log10_cal = 16'b0000010101110100;
            15'd23676: log10_cal = 16'b0000010101110100;
            15'd23677: log10_cal = 16'b0000010101110100;
            15'd23678: log10_cal = 16'b0000010101110100;
            15'd23679: log10_cal = 16'b0000010101110100;
            15'd23680: log10_cal = 16'b0000010101110100;
            15'd23681: log10_cal = 16'b0000010101110100;
            15'd23682: log10_cal = 16'b0000010101110100;
            15'd23683: log10_cal = 16'b0000010101110100;
            15'd23684: log10_cal = 16'b0000010101110100;
            15'd23685: log10_cal = 16'b0000010101110100;
            15'd23686: log10_cal = 16'b0000010101110100;
            15'd23687: log10_cal = 16'b0000010101110100;
            15'd23688: log10_cal = 16'b0000010101110100;
            15'd23689: log10_cal = 16'b0000010101110100;
            15'd23690: log10_cal = 16'b0000010101110101;
            15'd23691: log10_cal = 16'b0000010101110101;
            15'd23692: log10_cal = 16'b0000010101110101;
            15'd23693: log10_cal = 16'b0000010101110101;
            15'd23694: log10_cal = 16'b0000010101110101;
            15'd23695: log10_cal = 16'b0000010101110101;
            15'd23696: log10_cal = 16'b0000010101110101;
            15'd23697: log10_cal = 16'b0000010101110101;
            15'd23698: log10_cal = 16'b0000010101110101;
            15'd23699: log10_cal = 16'b0000010101110101;
            15'd23700: log10_cal = 16'b0000010101110101;
            15'd23701: log10_cal = 16'b0000010101110101;
            15'd23702: log10_cal = 16'b0000010101110101;
            15'd23703: log10_cal = 16'b0000010101110101;
            15'd23704: log10_cal = 16'b0000010101110101;
            15'd23705: log10_cal = 16'b0000010101110101;
            15'd23706: log10_cal = 16'b0000010101110101;
            15'd23707: log10_cal = 16'b0000010101110101;
            15'd23708: log10_cal = 16'b0000010101110101;
            15'd23709: log10_cal = 16'b0000010101110101;
            15'd23710: log10_cal = 16'b0000010101110101;
            15'd23711: log10_cal = 16'b0000010101110101;
            15'd23712: log10_cal = 16'b0000010101110101;
            15'd23713: log10_cal = 16'b0000010101110101;
            15'd23714: log10_cal = 16'b0000010101110101;
            15'd23715: log10_cal = 16'b0000010101110101;
            15'd23716: log10_cal = 16'b0000010101110101;
            15'd23717: log10_cal = 16'b0000010101110101;
            15'd23718: log10_cal = 16'b0000010101110101;
            15'd23719: log10_cal = 16'b0000010101110101;
            15'd23720: log10_cal = 16'b0000010101110101;
            15'd23721: log10_cal = 16'b0000010101110101;
            15'd23722: log10_cal = 16'b0000010101110101;
            15'd23723: log10_cal = 16'b0000010101110101;
            15'd23724: log10_cal = 16'b0000010101110101;
            15'd23725: log10_cal = 16'b0000010101110101;
            15'd23726: log10_cal = 16'b0000010101110101;
            15'd23727: log10_cal = 16'b0000010101110101;
            15'd23728: log10_cal = 16'b0000010101110101;
            15'd23729: log10_cal = 16'b0000010101110101;
            15'd23730: log10_cal = 16'b0000010101110101;
            15'd23731: log10_cal = 16'b0000010101110101;
            15'd23732: log10_cal = 16'b0000010101110101;
            15'd23733: log10_cal = 16'b0000010101110101;
            15'd23734: log10_cal = 16'b0000010101110101;
            15'd23735: log10_cal = 16'b0000010101110101;
            15'd23736: log10_cal = 16'b0000010101110101;
            15'd23737: log10_cal = 16'b0000010101110101;
            15'd23738: log10_cal = 16'b0000010101110101;
            15'd23739: log10_cal = 16'b0000010101110101;
            15'd23740: log10_cal = 16'b0000010101110101;
            15'd23741: log10_cal = 16'b0000010101110101;
            15'd23742: log10_cal = 16'b0000010101110101;
            15'd23743: log10_cal = 16'b0000010101110110;
            15'd23744: log10_cal = 16'b0000010101110110;
            15'd23745: log10_cal = 16'b0000010101110110;
            15'd23746: log10_cal = 16'b0000010101110110;
            15'd23747: log10_cal = 16'b0000010101110110;
            15'd23748: log10_cal = 16'b0000010101110110;
            15'd23749: log10_cal = 16'b0000010101110110;
            15'd23750: log10_cal = 16'b0000010101110110;
            15'd23751: log10_cal = 16'b0000010101110110;
            15'd23752: log10_cal = 16'b0000010101110110;
            15'd23753: log10_cal = 16'b0000010101110110;
            15'd23754: log10_cal = 16'b0000010101110110;
            15'd23755: log10_cal = 16'b0000010101110110;
            15'd23756: log10_cal = 16'b0000010101110110;
            15'd23757: log10_cal = 16'b0000010101110110;
            15'd23758: log10_cal = 16'b0000010101110110;
            15'd23759: log10_cal = 16'b0000010101110110;
            15'd23760: log10_cal = 16'b0000010101110110;
            15'd23761: log10_cal = 16'b0000010101110110;
            15'd23762: log10_cal = 16'b0000010101110110;
            15'd23763: log10_cal = 16'b0000010101110110;
            15'd23764: log10_cal = 16'b0000010101110110;
            15'd23765: log10_cal = 16'b0000010101110110;
            15'd23766: log10_cal = 16'b0000010101110110;
            15'd23767: log10_cal = 16'b0000010101110110;
            15'd23768: log10_cal = 16'b0000010101110110;
            15'd23769: log10_cal = 16'b0000010101110110;
            15'd23770: log10_cal = 16'b0000010101110110;
            15'd23771: log10_cal = 16'b0000010101110110;
            15'd23772: log10_cal = 16'b0000010101110110;
            15'd23773: log10_cal = 16'b0000010101110110;
            15'd23774: log10_cal = 16'b0000010101110110;
            15'd23775: log10_cal = 16'b0000010101110110;
            15'd23776: log10_cal = 16'b0000010101110110;
            15'd23777: log10_cal = 16'b0000010101110110;
            15'd23778: log10_cal = 16'b0000010101110110;
            15'd23779: log10_cal = 16'b0000010101110110;
            15'd23780: log10_cal = 16'b0000010101110110;
            15'd23781: log10_cal = 16'b0000010101110110;
            15'd23782: log10_cal = 16'b0000010101110110;
            15'd23783: log10_cal = 16'b0000010101110110;
            15'd23784: log10_cal = 16'b0000010101110110;
            15'd23785: log10_cal = 16'b0000010101110110;
            15'd23786: log10_cal = 16'b0000010101110110;
            15'd23787: log10_cal = 16'b0000010101110110;
            15'd23788: log10_cal = 16'b0000010101110110;
            15'd23789: log10_cal = 16'b0000010101110110;
            15'd23790: log10_cal = 16'b0000010101110110;
            15'd23791: log10_cal = 16'b0000010101110110;
            15'd23792: log10_cal = 16'b0000010101110110;
            15'd23793: log10_cal = 16'b0000010101110110;
            15'd23794: log10_cal = 16'b0000010101110110;
            15'd23795: log10_cal = 16'b0000010101110110;
            15'd23796: log10_cal = 16'b0000010101110110;
            15'd23797: log10_cal = 16'b0000010101110111;
            15'd23798: log10_cal = 16'b0000010101110111;
            15'd23799: log10_cal = 16'b0000010101110111;
            15'd23800: log10_cal = 16'b0000010101110111;
            15'd23801: log10_cal = 16'b0000010101110111;
            15'd23802: log10_cal = 16'b0000010101110111;
            15'd23803: log10_cal = 16'b0000010101110111;
            15'd23804: log10_cal = 16'b0000010101110111;
            15'd23805: log10_cal = 16'b0000010101110111;
            15'd23806: log10_cal = 16'b0000010101110111;
            15'd23807: log10_cal = 16'b0000010101110111;
            15'd23808: log10_cal = 16'b0000010101110111;
            15'd23809: log10_cal = 16'b0000010101110111;
            15'd23810: log10_cal = 16'b0000010101110111;
            15'd23811: log10_cal = 16'b0000010101110111;
            15'd23812: log10_cal = 16'b0000010101110111;
            15'd23813: log10_cal = 16'b0000010101110111;
            15'd23814: log10_cal = 16'b0000010101110111;
            15'd23815: log10_cal = 16'b0000010101110111;
            15'd23816: log10_cal = 16'b0000010101110111;
            15'd23817: log10_cal = 16'b0000010101110111;
            15'd23818: log10_cal = 16'b0000010101110111;
            15'd23819: log10_cal = 16'b0000010101110111;
            15'd23820: log10_cal = 16'b0000010101110111;
            15'd23821: log10_cal = 16'b0000010101110111;
            15'd23822: log10_cal = 16'b0000010101110111;
            15'd23823: log10_cal = 16'b0000010101110111;
            15'd23824: log10_cal = 16'b0000010101110111;
            15'd23825: log10_cal = 16'b0000010101110111;
            15'd23826: log10_cal = 16'b0000010101110111;
            15'd23827: log10_cal = 16'b0000010101110111;
            15'd23828: log10_cal = 16'b0000010101110111;
            15'd23829: log10_cal = 16'b0000010101110111;
            15'd23830: log10_cal = 16'b0000010101110111;
            15'd23831: log10_cal = 16'b0000010101110111;
            15'd23832: log10_cal = 16'b0000010101110111;
            15'd23833: log10_cal = 16'b0000010101110111;
            15'd23834: log10_cal = 16'b0000010101110111;
            15'd23835: log10_cal = 16'b0000010101110111;
            15'd23836: log10_cal = 16'b0000010101110111;
            15'd23837: log10_cal = 16'b0000010101110111;
            15'd23838: log10_cal = 16'b0000010101110111;
            15'd23839: log10_cal = 16'b0000010101110111;
            15'd23840: log10_cal = 16'b0000010101110111;
            15'd23841: log10_cal = 16'b0000010101110111;
            15'd23842: log10_cal = 16'b0000010101110111;
            15'd23843: log10_cal = 16'b0000010101110111;
            15'd23844: log10_cal = 16'b0000010101110111;
            15'd23845: log10_cal = 16'b0000010101110111;
            15'd23846: log10_cal = 16'b0000010101110111;
            15'd23847: log10_cal = 16'b0000010101110111;
            15'd23848: log10_cal = 16'b0000010101110111;
            15'd23849: log10_cal = 16'b0000010101110111;
            15'd23850: log10_cal = 16'b0000010101111000;
            15'd23851: log10_cal = 16'b0000010101111000;
            15'd23852: log10_cal = 16'b0000010101111000;
            15'd23853: log10_cal = 16'b0000010101111000;
            15'd23854: log10_cal = 16'b0000010101111000;
            15'd23855: log10_cal = 16'b0000010101111000;
            15'd23856: log10_cal = 16'b0000010101111000;
            15'd23857: log10_cal = 16'b0000010101111000;
            15'd23858: log10_cal = 16'b0000010101111000;
            15'd23859: log10_cal = 16'b0000010101111000;
            15'd23860: log10_cal = 16'b0000010101111000;
            15'd23861: log10_cal = 16'b0000010101111000;
            15'd23862: log10_cal = 16'b0000010101111000;
            15'd23863: log10_cal = 16'b0000010101111000;
            15'd23864: log10_cal = 16'b0000010101111000;
            15'd23865: log10_cal = 16'b0000010101111000;
            15'd23866: log10_cal = 16'b0000010101111000;
            15'd23867: log10_cal = 16'b0000010101111000;
            15'd23868: log10_cal = 16'b0000010101111000;
            15'd23869: log10_cal = 16'b0000010101111000;
            15'd23870: log10_cal = 16'b0000010101111000;
            15'd23871: log10_cal = 16'b0000010101111000;
            15'd23872: log10_cal = 16'b0000010101111000;
            15'd23873: log10_cal = 16'b0000010101111000;
            15'd23874: log10_cal = 16'b0000010101111000;
            15'd23875: log10_cal = 16'b0000010101111000;
            15'd23876: log10_cal = 16'b0000010101111000;
            15'd23877: log10_cal = 16'b0000010101111000;
            15'd23878: log10_cal = 16'b0000010101111000;
            15'd23879: log10_cal = 16'b0000010101111000;
            15'd23880: log10_cal = 16'b0000010101111000;
            15'd23881: log10_cal = 16'b0000010101111000;
            15'd23882: log10_cal = 16'b0000010101111000;
            15'd23883: log10_cal = 16'b0000010101111000;
            15'd23884: log10_cal = 16'b0000010101111000;
            15'd23885: log10_cal = 16'b0000010101111000;
            15'd23886: log10_cal = 16'b0000010101111000;
            15'd23887: log10_cal = 16'b0000010101111000;
            15'd23888: log10_cal = 16'b0000010101111000;
            15'd23889: log10_cal = 16'b0000010101111000;
            15'd23890: log10_cal = 16'b0000010101111000;
            15'd23891: log10_cal = 16'b0000010101111000;
            15'd23892: log10_cal = 16'b0000010101111000;
            15'd23893: log10_cal = 16'b0000010101111000;
            15'd23894: log10_cal = 16'b0000010101111000;
            15'd23895: log10_cal = 16'b0000010101111000;
            15'd23896: log10_cal = 16'b0000010101111000;
            15'd23897: log10_cal = 16'b0000010101111000;
            15'd23898: log10_cal = 16'b0000010101111000;
            15'd23899: log10_cal = 16'b0000010101111000;
            15'd23900: log10_cal = 16'b0000010101111000;
            15'd23901: log10_cal = 16'b0000010101111000;
            15'd23902: log10_cal = 16'b0000010101111000;
            15'd23903: log10_cal = 16'b0000010101111000;
            15'd23904: log10_cal = 16'b0000010101111001;
            15'd23905: log10_cal = 16'b0000010101111001;
            15'd23906: log10_cal = 16'b0000010101111001;
            15'd23907: log10_cal = 16'b0000010101111001;
            15'd23908: log10_cal = 16'b0000010101111001;
            15'd23909: log10_cal = 16'b0000010101111001;
            15'd23910: log10_cal = 16'b0000010101111001;
            15'd23911: log10_cal = 16'b0000010101111001;
            15'd23912: log10_cal = 16'b0000010101111001;
            15'd23913: log10_cal = 16'b0000010101111001;
            15'd23914: log10_cal = 16'b0000010101111001;
            15'd23915: log10_cal = 16'b0000010101111001;
            15'd23916: log10_cal = 16'b0000010101111001;
            15'd23917: log10_cal = 16'b0000010101111001;
            15'd23918: log10_cal = 16'b0000010101111001;
            15'd23919: log10_cal = 16'b0000010101111001;
            15'd23920: log10_cal = 16'b0000010101111001;
            15'd23921: log10_cal = 16'b0000010101111001;
            15'd23922: log10_cal = 16'b0000010101111001;
            15'd23923: log10_cal = 16'b0000010101111001;
            15'd23924: log10_cal = 16'b0000010101111001;
            15'd23925: log10_cal = 16'b0000010101111001;
            15'd23926: log10_cal = 16'b0000010101111001;
            15'd23927: log10_cal = 16'b0000010101111001;
            15'd23928: log10_cal = 16'b0000010101111001;
            15'd23929: log10_cal = 16'b0000010101111001;
            15'd23930: log10_cal = 16'b0000010101111001;
            15'd23931: log10_cal = 16'b0000010101111001;
            15'd23932: log10_cal = 16'b0000010101111001;
            15'd23933: log10_cal = 16'b0000010101111001;
            15'd23934: log10_cal = 16'b0000010101111001;
            15'd23935: log10_cal = 16'b0000010101111001;
            15'd23936: log10_cal = 16'b0000010101111001;
            15'd23937: log10_cal = 16'b0000010101111001;
            15'd23938: log10_cal = 16'b0000010101111001;
            15'd23939: log10_cal = 16'b0000010101111001;
            15'd23940: log10_cal = 16'b0000010101111001;
            15'd23941: log10_cal = 16'b0000010101111001;
            15'd23942: log10_cal = 16'b0000010101111001;
            15'd23943: log10_cal = 16'b0000010101111001;
            15'd23944: log10_cal = 16'b0000010101111001;
            15'd23945: log10_cal = 16'b0000010101111001;
            15'd23946: log10_cal = 16'b0000010101111001;
            15'd23947: log10_cal = 16'b0000010101111001;
            15'd23948: log10_cal = 16'b0000010101111001;
            15'd23949: log10_cal = 16'b0000010101111001;
            15'd23950: log10_cal = 16'b0000010101111001;
            15'd23951: log10_cal = 16'b0000010101111001;
            15'd23952: log10_cal = 16'b0000010101111001;
            15'd23953: log10_cal = 16'b0000010101111001;
            15'd23954: log10_cal = 16'b0000010101111001;
            15'd23955: log10_cal = 16'b0000010101111001;
            15'd23956: log10_cal = 16'b0000010101111001;
            15'd23957: log10_cal = 16'b0000010101111001;
            15'd23958: log10_cal = 16'b0000010101111010;
            15'd23959: log10_cal = 16'b0000010101111010;
            15'd23960: log10_cal = 16'b0000010101111010;
            15'd23961: log10_cal = 16'b0000010101111010;
            15'd23962: log10_cal = 16'b0000010101111010;
            15'd23963: log10_cal = 16'b0000010101111010;
            15'd23964: log10_cal = 16'b0000010101111010;
            15'd23965: log10_cal = 16'b0000010101111010;
            15'd23966: log10_cal = 16'b0000010101111010;
            15'd23967: log10_cal = 16'b0000010101111010;
            15'd23968: log10_cal = 16'b0000010101111010;
            15'd23969: log10_cal = 16'b0000010101111010;
            15'd23970: log10_cal = 16'b0000010101111010;
            15'd23971: log10_cal = 16'b0000010101111010;
            15'd23972: log10_cal = 16'b0000010101111010;
            15'd23973: log10_cal = 16'b0000010101111010;
            15'd23974: log10_cal = 16'b0000010101111010;
            15'd23975: log10_cal = 16'b0000010101111010;
            15'd23976: log10_cal = 16'b0000010101111010;
            15'd23977: log10_cal = 16'b0000010101111010;
            15'd23978: log10_cal = 16'b0000010101111010;
            15'd23979: log10_cal = 16'b0000010101111010;
            15'd23980: log10_cal = 16'b0000010101111010;
            15'd23981: log10_cal = 16'b0000010101111010;
            15'd23982: log10_cal = 16'b0000010101111010;
            15'd23983: log10_cal = 16'b0000010101111010;
            15'd23984: log10_cal = 16'b0000010101111010;
            15'd23985: log10_cal = 16'b0000010101111010;
            15'd23986: log10_cal = 16'b0000010101111010;
            15'd23987: log10_cal = 16'b0000010101111010;
            15'd23988: log10_cal = 16'b0000010101111010;
            15'd23989: log10_cal = 16'b0000010101111010;
            15'd23990: log10_cal = 16'b0000010101111010;
            15'd23991: log10_cal = 16'b0000010101111010;
            15'd23992: log10_cal = 16'b0000010101111010;
            15'd23993: log10_cal = 16'b0000010101111010;
            15'd23994: log10_cal = 16'b0000010101111010;
            15'd23995: log10_cal = 16'b0000010101111010;
            15'd23996: log10_cal = 16'b0000010101111010;
            15'd23997: log10_cal = 16'b0000010101111010;
            15'd23998: log10_cal = 16'b0000010101111010;
            15'd23999: log10_cal = 16'b0000010101111010;
            15'd24000: log10_cal = 16'b0000010101111010;
            15'd24001: log10_cal = 16'b0000010101111010;
            15'd24002: log10_cal = 16'b0000010101111010;
            15'd24003: log10_cal = 16'b0000010101111010;
            15'd24004: log10_cal = 16'b0000010101111010;
            15'd24005: log10_cal = 16'b0000010101111010;
            15'd24006: log10_cal = 16'b0000010101111010;
            15'd24007: log10_cal = 16'b0000010101111010;
            15'd24008: log10_cal = 16'b0000010101111010;
            15'd24009: log10_cal = 16'b0000010101111010;
            15'd24010: log10_cal = 16'b0000010101111010;
            15'd24011: log10_cal = 16'b0000010101111010;
            15'd24012: log10_cal = 16'b0000010101111011;
            15'd24013: log10_cal = 16'b0000010101111011;
            15'd24014: log10_cal = 16'b0000010101111011;
            15'd24015: log10_cal = 16'b0000010101111011;
            15'd24016: log10_cal = 16'b0000010101111011;
            15'd24017: log10_cal = 16'b0000010101111011;
            15'd24018: log10_cal = 16'b0000010101111011;
            15'd24019: log10_cal = 16'b0000010101111011;
            15'd24020: log10_cal = 16'b0000010101111011;
            15'd24021: log10_cal = 16'b0000010101111011;
            15'd24022: log10_cal = 16'b0000010101111011;
            15'd24023: log10_cal = 16'b0000010101111011;
            15'd24024: log10_cal = 16'b0000010101111011;
            15'd24025: log10_cal = 16'b0000010101111011;
            15'd24026: log10_cal = 16'b0000010101111011;
            15'd24027: log10_cal = 16'b0000010101111011;
            15'd24028: log10_cal = 16'b0000010101111011;
            15'd24029: log10_cal = 16'b0000010101111011;
            15'd24030: log10_cal = 16'b0000010101111011;
            15'd24031: log10_cal = 16'b0000010101111011;
            15'd24032: log10_cal = 16'b0000010101111011;
            15'd24033: log10_cal = 16'b0000010101111011;
            15'd24034: log10_cal = 16'b0000010101111011;
            15'd24035: log10_cal = 16'b0000010101111011;
            15'd24036: log10_cal = 16'b0000010101111011;
            15'd24037: log10_cal = 16'b0000010101111011;
            15'd24038: log10_cal = 16'b0000010101111011;
            15'd24039: log10_cal = 16'b0000010101111011;
            15'd24040: log10_cal = 16'b0000010101111011;
            15'd24041: log10_cal = 16'b0000010101111011;
            15'd24042: log10_cal = 16'b0000010101111011;
            15'd24043: log10_cal = 16'b0000010101111011;
            15'd24044: log10_cal = 16'b0000010101111011;
            15'd24045: log10_cal = 16'b0000010101111011;
            15'd24046: log10_cal = 16'b0000010101111011;
            15'd24047: log10_cal = 16'b0000010101111011;
            15'd24048: log10_cal = 16'b0000010101111011;
            15'd24049: log10_cal = 16'b0000010101111011;
            15'd24050: log10_cal = 16'b0000010101111011;
            15'd24051: log10_cal = 16'b0000010101111011;
            15'd24052: log10_cal = 16'b0000010101111011;
            15'd24053: log10_cal = 16'b0000010101111011;
            15'd24054: log10_cal = 16'b0000010101111011;
            15'd24055: log10_cal = 16'b0000010101111011;
            15'd24056: log10_cal = 16'b0000010101111011;
            15'd24057: log10_cal = 16'b0000010101111011;
            15'd24058: log10_cal = 16'b0000010101111011;
            15'd24059: log10_cal = 16'b0000010101111011;
            15'd24060: log10_cal = 16'b0000010101111011;
            15'd24061: log10_cal = 16'b0000010101111011;
            15'd24062: log10_cal = 16'b0000010101111011;
            15'd24063: log10_cal = 16'b0000010101111011;
            15'd24064: log10_cal = 16'b0000010101111011;
            15'd24065: log10_cal = 16'b0000010101111011;
            15'd24066: log10_cal = 16'b0000010101111100;
            15'd24067: log10_cal = 16'b0000010101111100;
            15'd24068: log10_cal = 16'b0000010101111100;
            15'd24069: log10_cal = 16'b0000010101111100;
            15'd24070: log10_cal = 16'b0000010101111100;
            15'd24071: log10_cal = 16'b0000010101111100;
            15'd24072: log10_cal = 16'b0000010101111100;
            15'd24073: log10_cal = 16'b0000010101111100;
            15'd24074: log10_cal = 16'b0000010101111100;
            15'd24075: log10_cal = 16'b0000010101111100;
            15'd24076: log10_cal = 16'b0000010101111100;
            15'd24077: log10_cal = 16'b0000010101111100;
            15'd24078: log10_cal = 16'b0000010101111100;
            15'd24079: log10_cal = 16'b0000010101111100;
            15'd24080: log10_cal = 16'b0000010101111100;
            15'd24081: log10_cal = 16'b0000010101111100;
            15'd24082: log10_cal = 16'b0000010101111100;
            15'd24083: log10_cal = 16'b0000010101111100;
            15'd24084: log10_cal = 16'b0000010101111100;
            15'd24085: log10_cal = 16'b0000010101111100;
            15'd24086: log10_cal = 16'b0000010101111100;
            15'd24087: log10_cal = 16'b0000010101111100;
            15'd24088: log10_cal = 16'b0000010101111100;
            15'd24089: log10_cal = 16'b0000010101111100;
            15'd24090: log10_cal = 16'b0000010101111100;
            15'd24091: log10_cal = 16'b0000010101111100;
            15'd24092: log10_cal = 16'b0000010101111100;
            15'd24093: log10_cal = 16'b0000010101111100;
            15'd24094: log10_cal = 16'b0000010101111100;
            15'd24095: log10_cal = 16'b0000010101111100;
            15'd24096: log10_cal = 16'b0000010101111100;
            15'd24097: log10_cal = 16'b0000010101111100;
            15'd24098: log10_cal = 16'b0000010101111100;
            15'd24099: log10_cal = 16'b0000010101111100;
            15'd24100: log10_cal = 16'b0000010101111100;
            15'd24101: log10_cal = 16'b0000010101111100;
            15'd24102: log10_cal = 16'b0000010101111100;
            15'd24103: log10_cal = 16'b0000010101111100;
            15'd24104: log10_cal = 16'b0000010101111100;
            15'd24105: log10_cal = 16'b0000010101111100;
            15'd24106: log10_cal = 16'b0000010101111100;
            15'd24107: log10_cal = 16'b0000010101111100;
            15'd24108: log10_cal = 16'b0000010101111100;
            15'd24109: log10_cal = 16'b0000010101111100;
            15'd24110: log10_cal = 16'b0000010101111100;
            15'd24111: log10_cal = 16'b0000010101111100;
            15'd24112: log10_cal = 16'b0000010101111100;
            15'd24113: log10_cal = 16'b0000010101111100;
            15'd24114: log10_cal = 16'b0000010101111100;
            15'd24115: log10_cal = 16'b0000010101111100;
            15'd24116: log10_cal = 16'b0000010101111100;
            15'd24117: log10_cal = 16'b0000010101111100;
            15'd24118: log10_cal = 16'b0000010101111100;
            15'd24119: log10_cal = 16'b0000010101111100;
            15'd24120: log10_cal = 16'b0000010101111101;
            15'd24121: log10_cal = 16'b0000010101111101;
            15'd24122: log10_cal = 16'b0000010101111101;
            15'd24123: log10_cal = 16'b0000010101111101;
            15'd24124: log10_cal = 16'b0000010101111101;
            15'd24125: log10_cal = 16'b0000010101111101;
            15'd24126: log10_cal = 16'b0000010101111101;
            15'd24127: log10_cal = 16'b0000010101111101;
            15'd24128: log10_cal = 16'b0000010101111101;
            15'd24129: log10_cal = 16'b0000010101111101;
            15'd24130: log10_cal = 16'b0000010101111101;
            15'd24131: log10_cal = 16'b0000010101111101;
            15'd24132: log10_cal = 16'b0000010101111101;
            15'd24133: log10_cal = 16'b0000010101111101;
            15'd24134: log10_cal = 16'b0000010101111101;
            15'd24135: log10_cal = 16'b0000010101111101;
            15'd24136: log10_cal = 16'b0000010101111101;
            15'd24137: log10_cal = 16'b0000010101111101;
            15'd24138: log10_cal = 16'b0000010101111101;
            15'd24139: log10_cal = 16'b0000010101111101;
            15'd24140: log10_cal = 16'b0000010101111101;
            15'd24141: log10_cal = 16'b0000010101111101;
            15'd24142: log10_cal = 16'b0000010101111101;
            15'd24143: log10_cal = 16'b0000010101111101;
            15'd24144: log10_cal = 16'b0000010101111101;
            15'd24145: log10_cal = 16'b0000010101111101;
            15'd24146: log10_cal = 16'b0000010101111101;
            15'd24147: log10_cal = 16'b0000010101111101;
            15'd24148: log10_cal = 16'b0000010101111101;
            15'd24149: log10_cal = 16'b0000010101111101;
            15'd24150: log10_cal = 16'b0000010101111101;
            15'd24151: log10_cal = 16'b0000010101111101;
            15'd24152: log10_cal = 16'b0000010101111101;
            15'd24153: log10_cal = 16'b0000010101111101;
            15'd24154: log10_cal = 16'b0000010101111101;
            15'd24155: log10_cal = 16'b0000010101111101;
            15'd24156: log10_cal = 16'b0000010101111101;
            15'd24157: log10_cal = 16'b0000010101111101;
            15'd24158: log10_cal = 16'b0000010101111101;
            15'd24159: log10_cal = 16'b0000010101111101;
            15'd24160: log10_cal = 16'b0000010101111101;
            15'd24161: log10_cal = 16'b0000010101111101;
            15'd24162: log10_cal = 16'b0000010101111101;
            15'd24163: log10_cal = 16'b0000010101111101;
            15'd24164: log10_cal = 16'b0000010101111101;
            15'd24165: log10_cal = 16'b0000010101111101;
            15'd24166: log10_cal = 16'b0000010101111101;
            15'd24167: log10_cal = 16'b0000010101111101;
            15'd24168: log10_cal = 16'b0000010101111101;
            15'd24169: log10_cal = 16'b0000010101111101;
            15'd24170: log10_cal = 16'b0000010101111101;
            15'd24171: log10_cal = 16'b0000010101111101;
            15'd24172: log10_cal = 16'b0000010101111101;
            15'd24173: log10_cal = 16'b0000010101111101;
            15'd24174: log10_cal = 16'b0000010101111110;
            15'd24175: log10_cal = 16'b0000010101111110;
            15'd24176: log10_cal = 16'b0000010101111110;
            15'd24177: log10_cal = 16'b0000010101111110;
            15'd24178: log10_cal = 16'b0000010101111110;
            15'd24179: log10_cal = 16'b0000010101111110;
            15'd24180: log10_cal = 16'b0000010101111110;
            15'd24181: log10_cal = 16'b0000010101111110;
            15'd24182: log10_cal = 16'b0000010101111110;
            15'd24183: log10_cal = 16'b0000010101111110;
            15'd24184: log10_cal = 16'b0000010101111110;
            15'd24185: log10_cal = 16'b0000010101111110;
            15'd24186: log10_cal = 16'b0000010101111110;
            15'd24187: log10_cal = 16'b0000010101111110;
            15'd24188: log10_cal = 16'b0000010101111110;
            15'd24189: log10_cal = 16'b0000010101111110;
            15'd24190: log10_cal = 16'b0000010101111110;
            15'd24191: log10_cal = 16'b0000010101111110;
            15'd24192: log10_cal = 16'b0000010101111110;
            15'd24193: log10_cal = 16'b0000010101111110;
            15'd24194: log10_cal = 16'b0000010101111110;
            15'd24195: log10_cal = 16'b0000010101111110;
            15'd24196: log10_cal = 16'b0000010101111110;
            15'd24197: log10_cal = 16'b0000010101111110;
            15'd24198: log10_cal = 16'b0000010101111110;
            15'd24199: log10_cal = 16'b0000010101111110;
            15'd24200: log10_cal = 16'b0000010101111110;
            15'd24201: log10_cal = 16'b0000010101111110;
            15'd24202: log10_cal = 16'b0000010101111110;
            15'd24203: log10_cal = 16'b0000010101111110;
            15'd24204: log10_cal = 16'b0000010101111110;
            15'd24205: log10_cal = 16'b0000010101111110;
            15'd24206: log10_cal = 16'b0000010101111110;
            15'd24207: log10_cal = 16'b0000010101111110;
            15'd24208: log10_cal = 16'b0000010101111110;
            15'd24209: log10_cal = 16'b0000010101111110;
            15'd24210: log10_cal = 16'b0000010101111110;
            15'd24211: log10_cal = 16'b0000010101111110;
            15'd24212: log10_cal = 16'b0000010101111110;
            15'd24213: log10_cal = 16'b0000010101111110;
            15'd24214: log10_cal = 16'b0000010101111110;
            15'd24215: log10_cal = 16'b0000010101111110;
            15'd24216: log10_cal = 16'b0000010101111110;
            15'd24217: log10_cal = 16'b0000010101111110;
            15'd24218: log10_cal = 16'b0000010101111110;
            15'd24219: log10_cal = 16'b0000010101111110;
            15'd24220: log10_cal = 16'b0000010101111110;
            15'd24221: log10_cal = 16'b0000010101111110;
            15'd24222: log10_cal = 16'b0000010101111110;
            15'd24223: log10_cal = 16'b0000010101111110;
            15'd24224: log10_cal = 16'b0000010101111110;
            15'd24225: log10_cal = 16'b0000010101111110;
            15'd24226: log10_cal = 16'b0000010101111110;
            15'd24227: log10_cal = 16'b0000010101111110;
            15'd24228: log10_cal = 16'b0000010101111110;
            15'd24229: log10_cal = 16'b0000010101111111;
            15'd24230: log10_cal = 16'b0000010101111111;
            15'd24231: log10_cal = 16'b0000010101111111;
            15'd24232: log10_cal = 16'b0000010101111111;
            15'd24233: log10_cal = 16'b0000010101111111;
            15'd24234: log10_cal = 16'b0000010101111111;
            15'd24235: log10_cal = 16'b0000010101111111;
            15'd24236: log10_cal = 16'b0000010101111111;
            15'd24237: log10_cal = 16'b0000010101111111;
            15'd24238: log10_cal = 16'b0000010101111111;
            15'd24239: log10_cal = 16'b0000010101111111;
            15'd24240: log10_cal = 16'b0000010101111111;
            15'd24241: log10_cal = 16'b0000010101111111;
            15'd24242: log10_cal = 16'b0000010101111111;
            15'd24243: log10_cal = 16'b0000010101111111;
            15'd24244: log10_cal = 16'b0000010101111111;
            15'd24245: log10_cal = 16'b0000010101111111;
            15'd24246: log10_cal = 16'b0000010101111111;
            15'd24247: log10_cal = 16'b0000010101111111;
            15'd24248: log10_cal = 16'b0000010101111111;
            15'd24249: log10_cal = 16'b0000010101111111;
            15'd24250: log10_cal = 16'b0000010101111111;
            15'd24251: log10_cal = 16'b0000010101111111;
            15'd24252: log10_cal = 16'b0000010101111111;
            15'd24253: log10_cal = 16'b0000010101111111;
            15'd24254: log10_cal = 16'b0000010101111111;
            15'd24255: log10_cal = 16'b0000010101111111;
            15'd24256: log10_cal = 16'b0000010101111111;
            15'd24257: log10_cal = 16'b0000010101111111;
            15'd24258: log10_cal = 16'b0000010101111111;
            15'd24259: log10_cal = 16'b0000010101111111;
            15'd24260: log10_cal = 16'b0000010101111111;
            15'd24261: log10_cal = 16'b0000010101111111;
            15'd24262: log10_cal = 16'b0000010101111111;
            15'd24263: log10_cal = 16'b0000010101111111;
            15'd24264: log10_cal = 16'b0000010101111111;
            15'd24265: log10_cal = 16'b0000010101111111;
            15'd24266: log10_cal = 16'b0000010101111111;
            15'd24267: log10_cal = 16'b0000010101111111;
            15'd24268: log10_cal = 16'b0000010101111111;
            15'd24269: log10_cal = 16'b0000010101111111;
            15'd24270: log10_cal = 16'b0000010101111111;
            15'd24271: log10_cal = 16'b0000010101111111;
            15'd24272: log10_cal = 16'b0000010101111111;
            15'd24273: log10_cal = 16'b0000010101111111;
            15'd24274: log10_cal = 16'b0000010101111111;
            15'd24275: log10_cal = 16'b0000010101111111;
            15'd24276: log10_cal = 16'b0000010101111111;
            15'd24277: log10_cal = 16'b0000010101111111;
            15'd24278: log10_cal = 16'b0000010101111111;
            15'd24279: log10_cal = 16'b0000010101111111;
            15'd24280: log10_cal = 16'b0000010101111111;
            15'd24281: log10_cal = 16'b0000010101111111;
            15'd24282: log10_cal = 16'b0000010101111111;
            15'd24283: log10_cal = 16'b0000010110000000;
            15'd24284: log10_cal = 16'b0000010110000000;
            15'd24285: log10_cal = 16'b0000010110000000;
            15'd24286: log10_cal = 16'b0000010110000000;
            15'd24287: log10_cal = 16'b0000010110000000;
            15'd24288: log10_cal = 16'b0000010110000000;
            15'd24289: log10_cal = 16'b0000010110000000;
            15'd24290: log10_cal = 16'b0000010110000000;
            15'd24291: log10_cal = 16'b0000010110000000;
            15'd24292: log10_cal = 16'b0000010110000000;
            15'd24293: log10_cal = 16'b0000010110000000;
            15'd24294: log10_cal = 16'b0000010110000000;
            15'd24295: log10_cal = 16'b0000010110000000;
            15'd24296: log10_cal = 16'b0000010110000000;
            15'd24297: log10_cal = 16'b0000010110000000;
            15'd24298: log10_cal = 16'b0000010110000000;
            15'd24299: log10_cal = 16'b0000010110000000;
            15'd24300: log10_cal = 16'b0000010110000000;
            15'd24301: log10_cal = 16'b0000010110000000;
            15'd24302: log10_cal = 16'b0000010110000000;
            15'd24303: log10_cal = 16'b0000010110000000;
            15'd24304: log10_cal = 16'b0000010110000000;
            15'd24305: log10_cal = 16'b0000010110000000;
            15'd24306: log10_cal = 16'b0000010110000000;
            15'd24307: log10_cal = 16'b0000010110000000;
            15'd24308: log10_cal = 16'b0000010110000000;
            15'd24309: log10_cal = 16'b0000010110000000;
            15'd24310: log10_cal = 16'b0000010110000000;
            15'd24311: log10_cal = 16'b0000010110000000;
            15'd24312: log10_cal = 16'b0000010110000000;
            15'd24313: log10_cal = 16'b0000010110000000;
            15'd24314: log10_cal = 16'b0000010110000000;
            15'd24315: log10_cal = 16'b0000010110000000;
            15'd24316: log10_cal = 16'b0000010110000000;
            15'd24317: log10_cal = 16'b0000010110000000;
            15'd24318: log10_cal = 16'b0000010110000000;
            15'd24319: log10_cal = 16'b0000010110000000;
            15'd24320: log10_cal = 16'b0000010110000000;
            15'd24321: log10_cal = 16'b0000010110000000;
            15'd24322: log10_cal = 16'b0000010110000000;
            15'd24323: log10_cal = 16'b0000010110000000;
            15'd24324: log10_cal = 16'b0000010110000000;
            15'd24325: log10_cal = 16'b0000010110000000;
            15'd24326: log10_cal = 16'b0000010110000000;
            15'd24327: log10_cal = 16'b0000010110000000;
            15'd24328: log10_cal = 16'b0000010110000000;
            15'd24329: log10_cal = 16'b0000010110000000;
            15'd24330: log10_cal = 16'b0000010110000000;
            15'd24331: log10_cal = 16'b0000010110000000;
            15'd24332: log10_cal = 16'b0000010110000000;
            15'd24333: log10_cal = 16'b0000010110000000;
            15'd24334: log10_cal = 16'b0000010110000000;
            15'd24335: log10_cal = 16'b0000010110000000;
            15'd24336: log10_cal = 16'b0000010110000000;
            15'd24337: log10_cal = 16'b0000010110000000;
            15'd24338: log10_cal = 16'b0000010110000001;
            15'd24339: log10_cal = 16'b0000010110000001;
            15'd24340: log10_cal = 16'b0000010110000001;
            15'd24341: log10_cal = 16'b0000010110000001;
            15'd24342: log10_cal = 16'b0000010110000001;
            15'd24343: log10_cal = 16'b0000010110000001;
            15'd24344: log10_cal = 16'b0000010110000001;
            15'd24345: log10_cal = 16'b0000010110000001;
            15'd24346: log10_cal = 16'b0000010110000001;
            15'd24347: log10_cal = 16'b0000010110000001;
            15'd24348: log10_cal = 16'b0000010110000001;
            15'd24349: log10_cal = 16'b0000010110000001;
            15'd24350: log10_cal = 16'b0000010110000001;
            15'd24351: log10_cal = 16'b0000010110000001;
            15'd24352: log10_cal = 16'b0000010110000001;
            15'd24353: log10_cal = 16'b0000010110000001;
            15'd24354: log10_cal = 16'b0000010110000001;
            15'd24355: log10_cal = 16'b0000010110000001;
            15'd24356: log10_cal = 16'b0000010110000001;
            15'd24357: log10_cal = 16'b0000010110000001;
            15'd24358: log10_cal = 16'b0000010110000001;
            15'd24359: log10_cal = 16'b0000010110000001;
            15'd24360: log10_cal = 16'b0000010110000001;
            15'd24361: log10_cal = 16'b0000010110000001;
            15'd24362: log10_cal = 16'b0000010110000001;
            15'd24363: log10_cal = 16'b0000010110000001;
            15'd24364: log10_cal = 16'b0000010110000001;
            15'd24365: log10_cal = 16'b0000010110000001;
            15'd24366: log10_cal = 16'b0000010110000001;
            15'd24367: log10_cal = 16'b0000010110000001;
            15'd24368: log10_cal = 16'b0000010110000001;
            15'd24369: log10_cal = 16'b0000010110000001;
            15'd24370: log10_cal = 16'b0000010110000001;
            15'd24371: log10_cal = 16'b0000010110000001;
            15'd24372: log10_cal = 16'b0000010110000001;
            15'd24373: log10_cal = 16'b0000010110000001;
            15'd24374: log10_cal = 16'b0000010110000001;
            15'd24375: log10_cal = 16'b0000010110000001;
            15'd24376: log10_cal = 16'b0000010110000001;
            15'd24377: log10_cal = 16'b0000010110000001;
            15'd24378: log10_cal = 16'b0000010110000001;
            15'd24379: log10_cal = 16'b0000010110000001;
            15'd24380: log10_cal = 16'b0000010110000001;
            15'd24381: log10_cal = 16'b0000010110000001;
            15'd24382: log10_cal = 16'b0000010110000001;
            15'd24383: log10_cal = 16'b0000010110000001;
            15'd24384: log10_cal = 16'b0000010110000001;
            15'd24385: log10_cal = 16'b0000010110000001;
            15'd24386: log10_cal = 16'b0000010110000001;
            15'd24387: log10_cal = 16'b0000010110000001;
            15'd24388: log10_cal = 16'b0000010110000001;
            15'd24389: log10_cal = 16'b0000010110000001;
            15'd24390: log10_cal = 16'b0000010110000001;
            15'd24391: log10_cal = 16'b0000010110000001;
            15'd24392: log10_cal = 16'b0000010110000001;
            15'd24393: log10_cal = 16'b0000010110000010;
            15'd24394: log10_cal = 16'b0000010110000010;
            15'd24395: log10_cal = 16'b0000010110000010;
            15'd24396: log10_cal = 16'b0000010110000010;
            15'd24397: log10_cal = 16'b0000010110000010;
            15'd24398: log10_cal = 16'b0000010110000010;
            15'd24399: log10_cal = 16'b0000010110000010;
            15'd24400: log10_cal = 16'b0000010110000010;
            15'd24401: log10_cal = 16'b0000010110000010;
            15'd24402: log10_cal = 16'b0000010110000010;
            15'd24403: log10_cal = 16'b0000010110000010;
            15'd24404: log10_cal = 16'b0000010110000010;
            15'd24405: log10_cal = 16'b0000010110000010;
            15'd24406: log10_cal = 16'b0000010110000010;
            15'd24407: log10_cal = 16'b0000010110000010;
            15'd24408: log10_cal = 16'b0000010110000010;
            15'd24409: log10_cal = 16'b0000010110000010;
            15'd24410: log10_cal = 16'b0000010110000010;
            15'd24411: log10_cal = 16'b0000010110000010;
            15'd24412: log10_cal = 16'b0000010110000010;
            15'd24413: log10_cal = 16'b0000010110000010;
            15'd24414: log10_cal = 16'b0000010110000010;
            15'd24415: log10_cal = 16'b0000010110000010;
            15'd24416: log10_cal = 16'b0000010110000010;
            15'd24417: log10_cal = 16'b0000010110000010;
            15'd24418: log10_cal = 16'b0000010110000010;
            15'd24419: log10_cal = 16'b0000010110000010;
            15'd24420: log10_cal = 16'b0000010110000010;
            15'd24421: log10_cal = 16'b0000010110000010;
            15'd24422: log10_cal = 16'b0000010110000010;
            15'd24423: log10_cal = 16'b0000010110000010;
            15'd24424: log10_cal = 16'b0000010110000010;
            15'd24425: log10_cal = 16'b0000010110000010;
            15'd24426: log10_cal = 16'b0000010110000010;
            15'd24427: log10_cal = 16'b0000010110000010;
            15'd24428: log10_cal = 16'b0000010110000010;
            15'd24429: log10_cal = 16'b0000010110000010;
            15'd24430: log10_cal = 16'b0000010110000010;
            15'd24431: log10_cal = 16'b0000010110000010;
            15'd24432: log10_cal = 16'b0000010110000010;
            15'd24433: log10_cal = 16'b0000010110000010;
            15'd24434: log10_cal = 16'b0000010110000010;
            15'd24435: log10_cal = 16'b0000010110000010;
            15'd24436: log10_cal = 16'b0000010110000010;
            15'd24437: log10_cal = 16'b0000010110000010;
            15'd24438: log10_cal = 16'b0000010110000010;
            15'd24439: log10_cal = 16'b0000010110000010;
            15'd24440: log10_cal = 16'b0000010110000010;
            15'd24441: log10_cal = 16'b0000010110000010;
            15'd24442: log10_cal = 16'b0000010110000010;
            15'd24443: log10_cal = 16'b0000010110000010;
            15'd24444: log10_cal = 16'b0000010110000010;
            15'd24445: log10_cal = 16'b0000010110000010;
            15'd24446: log10_cal = 16'b0000010110000010;
            15'd24447: log10_cal = 16'b0000010110000010;
            15'd24448: log10_cal = 16'b0000010110000011;
            15'd24449: log10_cal = 16'b0000010110000011;
            15'd24450: log10_cal = 16'b0000010110000011;
            15'd24451: log10_cal = 16'b0000010110000011;
            15'd24452: log10_cal = 16'b0000010110000011;
            15'd24453: log10_cal = 16'b0000010110000011;
            15'd24454: log10_cal = 16'b0000010110000011;
            15'd24455: log10_cal = 16'b0000010110000011;
            15'd24456: log10_cal = 16'b0000010110000011;
            15'd24457: log10_cal = 16'b0000010110000011;
            15'd24458: log10_cal = 16'b0000010110000011;
            15'd24459: log10_cal = 16'b0000010110000011;
            15'd24460: log10_cal = 16'b0000010110000011;
            15'd24461: log10_cal = 16'b0000010110000011;
            15'd24462: log10_cal = 16'b0000010110000011;
            15'd24463: log10_cal = 16'b0000010110000011;
            15'd24464: log10_cal = 16'b0000010110000011;
            15'd24465: log10_cal = 16'b0000010110000011;
            15'd24466: log10_cal = 16'b0000010110000011;
            15'd24467: log10_cal = 16'b0000010110000011;
            15'd24468: log10_cal = 16'b0000010110000011;
            15'd24469: log10_cal = 16'b0000010110000011;
            15'd24470: log10_cal = 16'b0000010110000011;
            15'd24471: log10_cal = 16'b0000010110000011;
            15'd24472: log10_cal = 16'b0000010110000011;
            15'd24473: log10_cal = 16'b0000010110000011;
            15'd24474: log10_cal = 16'b0000010110000011;
            15'd24475: log10_cal = 16'b0000010110000011;
            15'd24476: log10_cal = 16'b0000010110000011;
            15'd24477: log10_cal = 16'b0000010110000011;
            15'd24478: log10_cal = 16'b0000010110000011;
            15'd24479: log10_cal = 16'b0000010110000011;
            15'd24480: log10_cal = 16'b0000010110000011;
            15'd24481: log10_cal = 16'b0000010110000011;
            15'd24482: log10_cal = 16'b0000010110000011;
            15'd24483: log10_cal = 16'b0000010110000011;
            15'd24484: log10_cal = 16'b0000010110000011;
            15'd24485: log10_cal = 16'b0000010110000011;
            15'd24486: log10_cal = 16'b0000010110000011;
            15'd24487: log10_cal = 16'b0000010110000011;
            15'd24488: log10_cal = 16'b0000010110000011;
            15'd24489: log10_cal = 16'b0000010110000011;
            15'd24490: log10_cal = 16'b0000010110000011;
            15'd24491: log10_cal = 16'b0000010110000011;
            15'd24492: log10_cal = 16'b0000010110000011;
            15'd24493: log10_cal = 16'b0000010110000011;
            15'd24494: log10_cal = 16'b0000010110000011;
            15'd24495: log10_cal = 16'b0000010110000011;
            15'd24496: log10_cal = 16'b0000010110000011;
            15'd24497: log10_cal = 16'b0000010110000011;
            15'd24498: log10_cal = 16'b0000010110000011;
            15'd24499: log10_cal = 16'b0000010110000011;
            15'd24500: log10_cal = 16'b0000010110000011;
            15'd24501: log10_cal = 16'b0000010110000011;
            15'd24502: log10_cal = 16'b0000010110000011;
            15'd24503: log10_cal = 16'b0000010110000100;
            15'd24504: log10_cal = 16'b0000010110000100;
            15'd24505: log10_cal = 16'b0000010110000100;
            15'd24506: log10_cal = 16'b0000010110000100;
            15'd24507: log10_cal = 16'b0000010110000100;
            15'd24508: log10_cal = 16'b0000010110000100;
            15'd24509: log10_cal = 16'b0000010110000100;
            15'd24510: log10_cal = 16'b0000010110000100;
            15'd24511: log10_cal = 16'b0000010110000100;
            15'd24512: log10_cal = 16'b0000010110000100;
            15'd24513: log10_cal = 16'b0000010110000100;
            15'd24514: log10_cal = 16'b0000010110000100;
            15'd24515: log10_cal = 16'b0000010110000100;
            15'd24516: log10_cal = 16'b0000010110000100;
            15'd24517: log10_cal = 16'b0000010110000100;
            15'd24518: log10_cal = 16'b0000010110000100;
            15'd24519: log10_cal = 16'b0000010110000100;
            15'd24520: log10_cal = 16'b0000010110000100;
            15'd24521: log10_cal = 16'b0000010110000100;
            15'd24522: log10_cal = 16'b0000010110000100;
            15'd24523: log10_cal = 16'b0000010110000100;
            15'd24524: log10_cal = 16'b0000010110000100;
            15'd24525: log10_cal = 16'b0000010110000100;
            15'd24526: log10_cal = 16'b0000010110000100;
            15'd24527: log10_cal = 16'b0000010110000100;
            15'd24528: log10_cal = 16'b0000010110000100;
            15'd24529: log10_cal = 16'b0000010110000100;
            15'd24530: log10_cal = 16'b0000010110000100;
            15'd24531: log10_cal = 16'b0000010110000100;
            15'd24532: log10_cal = 16'b0000010110000100;
            15'd24533: log10_cal = 16'b0000010110000100;
            15'd24534: log10_cal = 16'b0000010110000100;
            15'd24535: log10_cal = 16'b0000010110000100;
            15'd24536: log10_cal = 16'b0000010110000100;
            15'd24537: log10_cal = 16'b0000010110000100;
            15'd24538: log10_cal = 16'b0000010110000100;
            15'd24539: log10_cal = 16'b0000010110000100;
            15'd24540: log10_cal = 16'b0000010110000100;
            15'd24541: log10_cal = 16'b0000010110000100;
            15'd24542: log10_cal = 16'b0000010110000100;
            15'd24543: log10_cal = 16'b0000010110000100;
            15'd24544: log10_cal = 16'b0000010110000100;
            15'd24545: log10_cal = 16'b0000010110000100;
            15'd24546: log10_cal = 16'b0000010110000100;
            15'd24547: log10_cal = 16'b0000010110000100;
            15'd24548: log10_cal = 16'b0000010110000100;
            15'd24549: log10_cal = 16'b0000010110000100;
            15'd24550: log10_cal = 16'b0000010110000100;
            15'd24551: log10_cal = 16'b0000010110000100;
            15'd24552: log10_cal = 16'b0000010110000100;
            15'd24553: log10_cal = 16'b0000010110000100;
            15'd24554: log10_cal = 16'b0000010110000100;
            15'd24555: log10_cal = 16'b0000010110000100;
            15'd24556: log10_cal = 16'b0000010110000100;
            15'd24557: log10_cal = 16'b0000010110000100;
            15'd24558: log10_cal = 16'b0000010110000101;
            15'd24559: log10_cal = 16'b0000010110000101;
            15'd24560: log10_cal = 16'b0000010110000101;
            15'd24561: log10_cal = 16'b0000010110000101;
            15'd24562: log10_cal = 16'b0000010110000101;
            15'd24563: log10_cal = 16'b0000010110000101;
            15'd24564: log10_cal = 16'b0000010110000101;
            15'd24565: log10_cal = 16'b0000010110000101;
            15'd24566: log10_cal = 16'b0000010110000101;
            15'd24567: log10_cal = 16'b0000010110000101;
            15'd24568: log10_cal = 16'b0000010110000101;
            15'd24569: log10_cal = 16'b0000010110000101;
            15'd24570: log10_cal = 16'b0000010110000101;
            15'd24571: log10_cal = 16'b0000010110000101;
            15'd24572: log10_cal = 16'b0000010110000101;
            15'd24573: log10_cal = 16'b0000010110000101;
            15'd24574: log10_cal = 16'b0000010110000101;
            15'd24575: log10_cal = 16'b0000010110000101;
            15'd24576: log10_cal = 16'b0000010110000101;
            15'd24577: log10_cal = 16'b0000010110000101;
            15'd24578: log10_cal = 16'b0000010110000101;
            15'd24579: log10_cal = 16'b0000010110000101;
            15'd24580: log10_cal = 16'b0000010110000101;
            15'd24581: log10_cal = 16'b0000010110000101;
            15'd24582: log10_cal = 16'b0000010110000101;
            15'd24583: log10_cal = 16'b0000010110000101;
            15'd24584: log10_cal = 16'b0000010110000101;
            15'd24585: log10_cal = 16'b0000010110000101;
            15'd24586: log10_cal = 16'b0000010110000101;
            15'd24587: log10_cal = 16'b0000010110000101;
            15'd24588: log10_cal = 16'b0000010110000101;
            15'd24589: log10_cal = 16'b0000010110000101;
            15'd24590: log10_cal = 16'b0000010110000101;
            15'd24591: log10_cal = 16'b0000010110000101;
            15'd24592: log10_cal = 16'b0000010110000101;
            15'd24593: log10_cal = 16'b0000010110000101;
            15'd24594: log10_cal = 16'b0000010110000101;
            15'd24595: log10_cal = 16'b0000010110000101;
            15'd24596: log10_cal = 16'b0000010110000101;
            15'd24597: log10_cal = 16'b0000010110000101;
            15'd24598: log10_cal = 16'b0000010110000101;
            15'd24599: log10_cal = 16'b0000010110000101;
            15'd24600: log10_cal = 16'b0000010110000101;
            15'd24601: log10_cal = 16'b0000010110000101;
            15'd24602: log10_cal = 16'b0000010110000101;
            15'd24603: log10_cal = 16'b0000010110000101;
            15'd24604: log10_cal = 16'b0000010110000101;
            15'd24605: log10_cal = 16'b0000010110000101;
            15'd24606: log10_cal = 16'b0000010110000101;
            15'd24607: log10_cal = 16'b0000010110000101;
            15'd24608: log10_cal = 16'b0000010110000101;
            15'd24609: log10_cal = 16'b0000010110000101;
            15'd24610: log10_cal = 16'b0000010110000101;
            15'd24611: log10_cal = 16'b0000010110000101;
            15'd24612: log10_cal = 16'b0000010110000101;
            15'd24613: log10_cal = 16'b0000010110000110;
            15'd24614: log10_cal = 16'b0000010110000110;
            15'd24615: log10_cal = 16'b0000010110000110;
            15'd24616: log10_cal = 16'b0000010110000110;
            15'd24617: log10_cal = 16'b0000010110000110;
            15'd24618: log10_cal = 16'b0000010110000110;
            15'd24619: log10_cal = 16'b0000010110000110;
            15'd24620: log10_cal = 16'b0000010110000110;
            15'd24621: log10_cal = 16'b0000010110000110;
            15'd24622: log10_cal = 16'b0000010110000110;
            15'd24623: log10_cal = 16'b0000010110000110;
            15'd24624: log10_cal = 16'b0000010110000110;
            15'd24625: log10_cal = 16'b0000010110000110;
            15'd24626: log10_cal = 16'b0000010110000110;
            15'd24627: log10_cal = 16'b0000010110000110;
            15'd24628: log10_cal = 16'b0000010110000110;
            15'd24629: log10_cal = 16'b0000010110000110;
            15'd24630: log10_cal = 16'b0000010110000110;
            15'd24631: log10_cal = 16'b0000010110000110;
            15'd24632: log10_cal = 16'b0000010110000110;
            15'd24633: log10_cal = 16'b0000010110000110;
            15'd24634: log10_cal = 16'b0000010110000110;
            15'd24635: log10_cal = 16'b0000010110000110;
            15'd24636: log10_cal = 16'b0000010110000110;
            15'd24637: log10_cal = 16'b0000010110000110;
            15'd24638: log10_cal = 16'b0000010110000110;
            15'd24639: log10_cal = 16'b0000010110000110;
            15'd24640: log10_cal = 16'b0000010110000110;
            15'd24641: log10_cal = 16'b0000010110000110;
            15'd24642: log10_cal = 16'b0000010110000110;
            15'd24643: log10_cal = 16'b0000010110000110;
            15'd24644: log10_cal = 16'b0000010110000110;
            15'd24645: log10_cal = 16'b0000010110000110;
            15'd24646: log10_cal = 16'b0000010110000110;
            15'd24647: log10_cal = 16'b0000010110000110;
            15'd24648: log10_cal = 16'b0000010110000110;
            15'd24649: log10_cal = 16'b0000010110000110;
            15'd24650: log10_cal = 16'b0000010110000110;
            15'd24651: log10_cal = 16'b0000010110000110;
            15'd24652: log10_cal = 16'b0000010110000110;
            15'd24653: log10_cal = 16'b0000010110000110;
            15'd24654: log10_cal = 16'b0000010110000110;
            15'd24655: log10_cal = 16'b0000010110000110;
            15'd24656: log10_cal = 16'b0000010110000110;
            15'd24657: log10_cal = 16'b0000010110000110;
            15'd24658: log10_cal = 16'b0000010110000110;
            15'd24659: log10_cal = 16'b0000010110000110;
            15'd24660: log10_cal = 16'b0000010110000110;
            15'd24661: log10_cal = 16'b0000010110000110;
            15'd24662: log10_cal = 16'b0000010110000110;
            15'd24663: log10_cal = 16'b0000010110000110;
            15'd24664: log10_cal = 16'b0000010110000110;
            15'd24665: log10_cal = 16'b0000010110000110;
            15'd24666: log10_cal = 16'b0000010110000110;
            15'd24667: log10_cal = 16'b0000010110000110;
            15'd24668: log10_cal = 16'b0000010110000110;
            15'd24669: log10_cal = 16'b0000010110000111;
            15'd24670: log10_cal = 16'b0000010110000111;
            15'd24671: log10_cal = 16'b0000010110000111;
            15'd24672: log10_cal = 16'b0000010110000111;
            15'd24673: log10_cal = 16'b0000010110000111;
            15'd24674: log10_cal = 16'b0000010110000111;
            15'd24675: log10_cal = 16'b0000010110000111;
            15'd24676: log10_cal = 16'b0000010110000111;
            15'd24677: log10_cal = 16'b0000010110000111;
            15'd24678: log10_cal = 16'b0000010110000111;
            15'd24679: log10_cal = 16'b0000010110000111;
            15'd24680: log10_cal = 16'b0000010110000111;
            15'd24681: log10_cal = 16'b0000010110000111;
            15'd24682: log10_cal = 16'b0000010110000111;
            15'd24683: log10_cal = 16'b0000010110000111;
            15'd24684: log10_cal = 16'b0000010110000111;
            15'd24685: log10_cal = 16'b0000010110000111;
            15'd24686: log10_cal = 16'b0000010110000111;
            15'd24687: log10_cal = 16'b0000010110000111;
            15'd24688: log10_cal = 16'b0000010110000111;
            15'd24689: log10_cal = 16'b0000010110000111;
            15'd24690: log10_cal = 16'b0000010110000111;
            15'd24691: log10_cal = 16'b0000010110000111;
            15'd24692: log10_cal = 16'b0000010110000111;
            15'd24693: log10_cal = 16'b0000010110000111;
            15'd24694: log10_cal = 16'b0000010110000111;
            15'd24695: log10_cal = 16'b0000010110000111;
            15'd24696: log10_cal = 16'b0000010110000111;
            15'd24697: log10_cal = 16'b0000010110000111;
            15'd24698: log10_cal = 16'b0000010110000111;
            15'd24699: log10_cal = 16'b0000010110000111;
            15'd24700: log10_cal = 16'b0000010110000111;
            15'd24701: log10_cal = 16'b0000010110000111;
            15'd24702: log10_cal = 16'b0000010110000111;
            15'd24703: log10_cal = 16'b0000010110000111;
            15'd24704: log10_cal = 16'b0000010110000111;
            15'd24705: log10_cal = 16'b0000010110000111;
            15'd24706: log10_cal = 16'b0000010110000111;
            15'd24707: log10_cal = 16'b0000010110000111;
            15'd24708: log10_cal = 16'b0000010110000111;
            15'd24709: log10_cal = 16'b0000010110000111;
            15'd24710: log10_cal = 16'b0000010110000111;
            15'd24711: log10_cal = 16'b0000010110000111;
            15'd24712: log10_cal = 16'b0000010110000111;
            15'd24713: log10_cal = 16'b0000010110000111;
            15'd24714: log10_cal = 16'b0000010110000111;
            15'd24715: log10_cal = 16'b0000010110000111;
            15'd24716: log10_cal = 16'b0000010110000111;
            15'd24717: log10_cal = 16'b0000010110000111;
            15'd24718: log10_cal = 16'b0000010110000111;
            15'd24719: log10_cal = 16'b0000010110000111;
            15'd24720: log10_cal = 16'b0000010110000111;
            15'd24721: log10_cal = 16'b0000010110000111;
            15'd24722: log10_cal = 16'b0000010110000111;
            15'd24723: log10_cal = 16'b0000010110000111;
            15'd24724: log10_cal = 16'b0000010110001000;
            15'd24725: log10_cal = 16'b0000010110001000;
            15'd24726: log10_cal = 16'b0000010110001000;
            15'd24727: log10_cal = 16'b0000010110001000;
            15'd24728: log10_cal = 16'b0000010110001000;
            15'd24729: log10_cal = 16'b0000010110001000;
            15'd24730: log10_cal = 16'b0000010110001000;
            15'd24731: log10_cal = 16'b0000010110001000;
            15'd24732: log10_cal = 16'b0000010110001000;
            15'd24733: log10_cal = 16'b0000010110001000;
            15'd24734: log10_cal = 16'b0000010110001000;
            15'd24735: log10_cal = 16'b0000010110001000;
            15'd24736: log10_cal = 16'b0000010110001000;
            15'd24737: log10_cal = 16'b0000010110001000;
            15'd24738: log10_cal = 16'b0000010110001000;
            15'd24739: log10_cal = 16'b0000010110001000;
            15'd24740: log10_cal = 16'b0000010110001000;
            15'd24741: log10_cal = 16'b0000010110001000;
            15'd24742: log10_cal = 16'b0000010110001000;
            15'd24743: log10_cal = 16'b0000010110001000;
            15'd24744: log10_cal = 16'b0000010110001000;
            15'd24745: log10_cal = 16'b0000010110001000;
            15'd24746: log10_cal = 16'b0000010110001000;
            15'd24747: log10_cal = 16'b0000010110001000;
            15'd24748: log10_cal = 16'b0000010110001000;
            15'd24749: log10_cal = 16'b0000010110001000;
            15'd24750: log10_cal = 16'b0000010110001000;
            15'd24751: log10_cal = 16'b0000010110001000;
            15'd24752: log10_cal = 16'b0000010110001000;
            15'd24753: log10_cal = 16'b0000010110001000;
            15'd24754: log10_cal = 16'b0000010110001000;
            15'd24755: log10_cal = 16'b0000010110001000;
            15'd24756: log10_cal = 16'b0000010110001000;
            15'd24757: log10_cal = 16'b0000010110001000;
            15'd24758: log10_cal = 16'b0000010110001000;
            15'd24759: log10_cal = 16'b0000010110001000;
            15'd24760: log10_cal = 16'b0000010110001000;
            15'd24761: log10_cal = 16'b0000010110001000;
            15'd24762: log10_cal = 16'b0000010110001000;
            15'd24763: log10_cal = 16'b0000010110001000;
            15'd24764: log10_cal = 16'b0000010110001000;
            15'd24765: log10_cal = 16'b0000010110001000;
            15'd24766: log10_cal = 16'b0000010110001000;
            15'd24767: log10_cal = 16'b0000010110001000;
            15'd24768: log10_cal = 16'b0000010110001000;
            15'd24769: log10_cal = 16'b0000010110001000;
            15'd24770: log10_cal = 16'b0000010110001000;
            15'd24771: log10_cal = 16'b0000010110001000;
            15'd24772: log10_cal = 16'b0000010110001000;
            15'd24773: log10_cal = 16'b0000010110001000;
            15'd24774: log10_cal = 16'b0000010110001000;
            15'd24775: log10_cal = 16'b0000010110001000;
            15'd24776: log10_cal = 16'b0000010110001000;
            15'd24777: log10_cal = 16'b0000010110001000;
            15'd24778: log10_cal = 16'b0000010110001000;
            15'd24779: log10_cal = 16'b0000010110001000;
            15'd24780: log10_cal = 16'b0000010110001001;
            15'd24781: log10_cal = 16'b0000010110001001;
            15'd24782: log10_cal = 16'b0000010110001001;
            15'd24783: log10_cal = 16'b0000010110001001;
            15'd24784: log10_cal = 16'b0000010110001001;
            15'd24785: log10_cal = 16'b0000010110001001;
            15'd24786: log10_cal = 16'b0000010110001001;
            15'd24787: log10_cal = 16'b0000010110001001;
            15'd24788: log10_cal = 16'b0000010110001001;
            15'd24789: log10_cal = 16'b0000010110001001;
            15'd24790: log10_cal = 16'b0000010110001001;
            15'd24791: log10_cal = 16'b0000010110001001;
            15'd24792: log10_cal = 16'b0000010110001001;
            15'd24793: log10_cal = 16'b0000010110001001;
            15'd24794: log10_cal = 16'b0000010110001001;
            15'd24795: log10_cal = 16'b0000010110001001;
            15'd24796: log10_cal = 16'b0000010110001001;
            15'd24797: log10_cal = 16'b0000010110001001;
            15'd24798: log10_cal = 16'b0000010110001001;
            15'd24799: log10_cal = 16'b0000010110001001;
            15'd24800: log10_cal = 16'b0000010110001001;
            15'd24801: log10_cal = 16'b0000010110001001;
            15'd24802: log10_cal = 16'b0000010110001001;
            15'd24803: log10_cal = 16'b0000010110001001;
            15'd24804: log10_cal = 16'b0000010110001001;
            15'd24805: log10_cal = 16'b0000010110001001;
            15'd24806: log10_cal = 16'b0000010110001001;
            15'd24807: log10_cal = 16'b0000010110001001;
            15'd24808: log10_cal = 16'b0000010110001001;
            15'd24809: log10_cal = 16'b0000010110001001;
            15'd24810: log10_cal = 16'b0000010110001001;
            15'd24811: log10_cal = 16'b0000010110001001;
            15'd24812: log10_cal = 16'b0000010110001001;
            15'd24813: log10_cal = 16'b0000010110001001;
            15'd24814: log10_cal = 16'b0000010110001001;
            15'd24815: log10_cal = 16'b0000010110001001;
            15'd24816: log10_cal = 16'b0000010110001001;
            15'd24817: log10_cal = 16'b0000010110001001;
            15'd24818: log10_cal = 16'b0000010110001001;
            15'd24819: log10_cal = 16'b0000010110001001;
            15'd24820: log10_cal = 16'b0000010110001001;
            15'd24821: log10_cal = 16'b0000010110001001;
            15'd24822: log10_cal = 16'b0000010110001001;
            15'd24823: log10_cal = 16'b0000010110001001;
            15'd24824: log10_cal = 16'b0000010110001001;
            15'd24825: log10_cal = 16'b0000010110001001;
            15'd24826: log10_cal = 16'b0000010110001001;
            15'd24827: log10_cal = 16'b0000010110001001;
            15'd24828: log10_cal = 16'b0000010110001001;
            15'd24829: log10_cal = 16'b0000010110001001;
            15'd24830: log10_cal = 16'b0000010110001001;
            15'd24831: log10_cal = 16'b0000010110001001;
            15'd24832: log10_cal = 16'b0000010110001001;
            15'd24833: log10_cal = 16'b0000010110001001;
            15'd24834: log10_cal = 16'b0000010110001001;
            15'd24835: log10_cal = 16'b0000010110001001;
            15'd24836: log10_cal = 16'b0000010110001010;
            15'd24837: log10_cal = 16'b0000010110001010;
            15'd24838: log10_cal = 16'b0000010110001010;
            15'd24839: log10_cal = 16'b0000010110001010;
            15'd24840: log10_cal = 16'b0000010110001010;
            15'd24841: log10_cal = 16'b0000010110001010;
            15'd24842: log10_cal = 16'b0000010110001010;
            15'd24843: log10_cal = 16'b0000010110001010;
            15'd24844: log10_cal = 16'b0000010110001010;
            15'd24845: log10_cal = 16'b0000010110001010;
            15'd24846: log10_cal = 16'b0000010110001010;
            15'd24847: log10_cal = 16'b0000010110001010;
            15'd24848: log10_cal = 16'b0000010110001010;
            15'd24849: log10_cal = 16'b0000010110001010;
            15'd24850: log10_cal = 16'b0000010110001010;
            15'd24851: log10_cal = 16'b0000010110001010;
            15'd24852: log10_cal = 16'b0000010110001010;
            15'd24853: log10_cal = 16'b0000010110001010;
            15'd24854: log10_cal = 16'b0000010110001010;
            15'd24855: log10_cal = 16'b0000010110001010;
            15'd24856: log10_cal = 16'b0000010110001010;
            15'd24857: log10_cal = 16'b0000010110001010;
            15'd24858: log10_cal = 16'b0000010110001010;
            15'd24859: log10_cal = 16'b0000010110001010;
            15'd24860: log10_cal = 16'b0000010110001010;
            15'd24861: log10_cal = 16'b0000010110001010;
            15'd24862: log10_cal = 16'b0000010110001010;
            15'd24863: log10_cal = 16'b0000010110001010;
            15'd24864: log10_cal = 16'b0000010110001010;
            15'd24865: log10_cal = 16'b0000010110001010;
            15'd24866: log10_cal = 16'b0000010110001010;
            15'd24867: log10_cal = 16'b0000010110001010;
            15'd24868: log10_cal = 16'b0000010110001010;
            15'd24869: log10_cal = 16'b0000010110001010;
            15'd24870: log10_cal = 16'b0000010110001010;
            15'd24871: log10_cal = 16'b0000010110001010;
            15'd24872: log10_cal = 16'b0000010110001010;
            15'd24873: log10_cal = 16'b0000010110001010;
            15'd24874: log10_cal = 16'b0000010110001010;
            15'd24875: log10_cal = 16'b0000010110001010;
            15'd24876: log10_cal = 16'b0000010110001010;
            15'd24877: log10_cal = 16'b0000010110001010;
            15'd24878: log10_cal = 16'b0000010110001010;
            15'd24879: log10_cal = 16'b0000010110001010;
            15'd24880: log10_cal = 16'b0000010110001010;
            15'd24881: log10_cal = 16'b0000010110001010;
            15'd24882: log10_cal = 16'b0000010110001010;
            15'd24883: log10_cal = 16'b0000010110001010;
            15'd24884: log10_cal = 16'b0000010110001010;
            15'd24885: log10_cal = 16'b0000010110001010;
            15'd24886: log10_cal = 16'b0000010110001010;
            15'd24887: log10_cal = 16'b0000010110001010;
            15'd24888: log10_cal = 16'b0000010110001010;
            15'd24889: log10_cal = 16'b0000010110001010;
            15'd24890: log10_cal = 16'b0000010110001010;
            15'd24891: log10_cal = 16'b0000010110001011;
            15'd24892: log10_cal = 16'b0000010110001011;
            15'd24893: log10_cal = 16'b0000010110001011;
            15'd24894: log10_cal = 16'b0000010110001011;
            15'd24895: log10_cal = 16'b0000010110001011;
            15'd24896: log10_cal = 16'b0000010110001011;
            15'd24897: log10_cal = 16'b0000010110001011;
            15'd24898: log10_cal = 16'b0000010110001011;
            15'd24899: log10_cal = 16'b0000010110001011;
            15'd24900: log10_cal = 16'b0000010110001011;
            15'd24901: log10_cal = 16'b0000010110001011;
            15'd24902: log10_cal = 16'b0000010110001011;
            15'd24903: log10_cal = 16'b0000010110001011;
            15'd24904: log10_cal = 16'b0000010110001011;
            15'd24905: log10_cal = 16'b0000010110001011;
            15'd24906: log10_cal = 16'b0000010110001011;
            15'd24907: log10_cal = 16'b0000010110001011;
            15'd24908: log10_cal = 16'b0000010110001011;
            15'd24909: log10_cal = 16'b0000010110001011;
            15'd24910: log10_cal = 16'b0000010110001011;
            15'd24911: log10_cal = 16'b0000010110001011;
            15'd24912: log10_cal = 16'b0000010110001011;
            15'd24913: log10_cal = 16'b0000010110001011;
            15'd24914: log10_cal = 16'b0000010110001011;
            15'd24915: log10_cal = 16'b0000010110001011;
            15'd24916: log10_cal = 16'b0000010110001011;
            15'd24917: log10_cal = 16'b0000010110001011;
            15'd24918: log10_cal = 16'b0000010110001011;
            15'd24919: log10_cal = 16'b0000010110001011;
            15'd24920: log10_cal = 16'b0000010110001011;
            15'd24921: log10_cal = 16'b0000010110001011;
            15'd24922: log10_cal = 16'b0000010110001011;
            15'd24923: log10_cal = 16'b0000010110001011;
            15'd24924: log10_cal = 16'b0000010110001011;
            15'd24925: log10_cal = 16'b0000010110001011;
            15'd24926: log10_cal = 16'b0000010110001011;
            15'd24927: log10_cal = 16'b0000010110001011;
            15'd24928: log10_cal = 16'b0000010110001011;
            15'd24929: log10_cal = 16'b0000010110001011;
            15'd24930: log10_cal = 16'b0000010110001011;
            15'd24931: log10_cal = 16'b0000010110001011;
            15'd24932: log10_cal = 16'b0000010110001011;
            15'd24933: log10_cal = 16'b0000010110001011;
            15'd24934: log10_cal = 16'b0000010110001011;
            15'd24935: log10_cal = 16'b0000010110001011;
            15'd24936: log10_cal = 16'b0000010110001011;
            15'd24937: log10_cal = 16'b0000010110001011;
            15'd24938: log10_cal = 16'b0000010110001011;
            15'd24939: log10_cal = 16'b0000010110001011;
            15'd24940: log10_cal = 16'b0000010110001011;
            15'd24941: log10_cal = 16'b0000010110001011;
            15'd24942: log10_cal = 16'b0000010110001011;
            15'd24943: log10_cal = 16'b0000010110001011;
            15'd24944: log10_cal = 16'b0000010110001011;
            15'd24945: log10_cal = 16'b0000010110001011;
            15'd24946: log10_cal = 16'b0000010110001011;
            15'd24947: log10_cal = 16'b0000010110001011;
            15'd24948: log10_cal = 16'b0000010110001100;
            15'd24949: log10_cal = 16'b0000010110001100;
            15'd24950: log10_cal = 16'b0000010110001100;
            15'd24951: log10_cal = 16'b0000010110001100;
            15'd24952: log10_cal = 16'b0000010110001100;
            15'd24953: log10_cal = 16'b0000010110001100;
            15'd24954: log10_cal = 16'b0000010110001100;
            15'd24955: log10_cal = 16'b0000010110001100;
            15'd24956: log10_cal = 16'b0000010110001100;
            15'd24957: log10_cal = 16'b0000010110001100;
            15'd24958: log10_cal = 16'b0000010110001100;
            15'd24959: log10_cal = 16'b0000010110001100;
            15'd24960: log10_cal = 16'b0000010110001100;
            15'd24961: log10_cal = 16'b0000010110001100;
            15'd24962: log10_cal = 16'b0000010110001100;
            15'd24963: log10_cal = 16'b0000010110001100;
            15'd24964: log10_cal = 16'b0000010110001100;
            15'd24965: log10_cal = 16'b0000010110001100;
            15'd24966: log10_cal = 16'b0000010110001100;
            15'd24967: log10_cal = 16'b0000010110001100;
            15'd24968: log10_cal = 16'b0000010110001100;
            15'd24969: log10_cal = 16'b0000010110001100;
            15'd24970: log10_cal = 16'b0000010110001100;
            15'd24971: log10_cal = 16'b0000010110001100;
            15'd24972: log10_cal = 16'b0000010110001100;
            15'd24973: log10_cal = 16'b0000010110001100;
            15'd24974: log10_cal = 16'b0000010110001100;
            15'd24975: log10_cal = 16'b0000010110001100;
            15'd24976: log10_cal = 16'b0000010110001100;
            15'd24977: log10_cal = 16'b0000010110001100;
            15'd24978: log10_cal = 16'b0000010110001100;
            15'd24979: log10_cal = 16'b0000010110001100;
            15'd24980: log10_cal = 16'b0000010110001100;
            15'd24981: log10_cal = 16'b0000010110001100;
            15'd24982: log10_cal = 16'b0000010110001100;
            15'd24983: log10_cal = 16'b0000010110001100;
            15'd24984: log10_cal = 16'b0000010110001100;
            15'd24985: log10_cal = 16'b0000010110001100;
            15'd24986: log10_cal = 16'b0000010110001100;
            15'd24987: log10_cal = 16'b0000010110001100;
            15'd24988: log10_cal = 16'b0000010110001100;
            15'd24989: log10_cal = 16'b0000010110001100;
            15'd24990: log10_cal = 16'b0000010110001100;
            15'd24991: log10_cal = 16'b0000010110001100;
            15'd24992: log10_cal = 16'b0000010110001100;
            15'd24993: log10_cal = 16'b0000010110001100;
            15'd24994: log10_cal = 16'b0000010110001100;
            15'd24995: log10_cal = 16'b0000010110001100;
            15'd24996: log10_cal = 16'b0000010110001100;
            15'd24997: log10_cal = 16'b0000010110001100;
            15'd24998: log10_cal = 16'b0000010110001100;
            15'd24999: log10_cal = 16'b0000010110001100;
            15'd25000: log10_cal = 16'b0000010110001100;
            15'd25001: log10_cal = 16'b0000010110001100;
            15'd25002: log10_cal = 16'b0000010110001100;
            15'd25003: log10_cal = 16'b0000010110001100;
            15'd25004: log10_cal = 16'b0000010110001101;
            15'd25005: log10_cal = 16'b0000010110001101;
            15'd25006: log10_cal = 16'b0000010110001101;
            15'd25007: log10_cal = 16'b0000010110001101;
            15'd25008: log10_cal = 16'b0000010110001101;
            15'd25009: log10_cal = 16'b0000010110001101;
            15'd25010: log10_cal = 16'b0000010110001101;
            15'd25011: log10_cal = 16'b0000010110001101;
            15'd25012: log10_cal = 16'b0000010110001101;
            15'd25013: log10_cal = 16'b0000010110001101;
            15'd25014: log10_cal = 16'b0000010110001101;
            15'd25015: log10_cal = 16'b0000010110001101;
            15'd25016: log10_cal = 16'b0000010110001101;
            15'd25017: log10_cal = 16'b0000010110001101;
            15'd25018: log10_cal = 16'b0000010110001101;
            15'd25019: log10_cal = 16'b0000010110001101;
            15'd25020: log10_cal = 16'b0000010110001101;
            15'd25021: log10_cal = 16'b0000010110001101;
            15'd25022: log10_cal = 16'b0000010110001101;
            15'd25023: log10_cal = 16'b0000010110001101;
            15'd25024: log10_cal = 16'b0000010110001101;
            15'd25025: log10_cal = 16'b0000010110001101;
            15'd25026: log10_cal = 16'b0000010110001101;
            15'd25027: log10_cal = 16'b0000010110001101;
            15'd25028: log10_cal = 16'b0000010110001101;
            15'd25029: log10_cal = 16'b0000010110001101;
            15'd25030: log10_cal = 16'b0000010110001101;
            15'd25031: log10_cal = 16'b0000010110001101;
            15'd25032: log10_cal = 16'b0000010110001101;
            15'd25033: log10_cal = 16'b0000010110001101;
            15'd25034: log10_cal = 16'b0000010110001101;
            15'd25035: log10_cal = 16'b0000010110001101;
            15'd25036: log10_cal = 16'b0000010110001101;
            15'd25037: log10_cal = 16'b0000010110001101;
            15'd25038: log10_cal = 16'b0000010110001101;
            15'd25039: log10_cal = 16'b0000010110001101;
            15'd25040: log10_cal = 16'b0000010110001101;
            15'd25041: log10_cal = 16'b0000010110001101;
            15'd25042: log10_cal = 16'b0000010110001101;
            15'd25043: log10_cal = 16'b0000010110001101;
            15'd25044: log10_cal = 16'b0000010110001101;
            15'd25045: log10_cal = 16'b0000010110001101;
            15'd25046: log10_cal = 16'b0000010110001101;
            15'd25047: log10_cal = 16'b0000010110001101;
            15'd25048: log10_cal = 16'b0000010110001101;
            15'd25049: log10_cal = 16'b0000010110001101;
            15'd25050: log10_cal = 16'b0000010110001101;
            15'd25051: log10_cal = 16'b0000010110001101;
            15'd25052: log10_cal = 16'b0000010110001101;
            15'd25053: log10_cal = 16'b0000010110001101;
            15'd25054: log10_cal = 16'b0000010110001101;
            15'd25055: log10_cal = 16'b0000010110001101;
            15'd25056: log10_cal = 16'b0000010110001101;
            15'd25057: log10_cal = 16'b0000010110001101;
            15'd25058: log10_cal = 16'b0000010110001101;
            15'd25059: log10_cal = 16'b0000010110001101;
            15'd25060: log10_cal = 16'b0000010110001110;
            15'd25061: log10_cal = 16'b0000010110001110;
            15'd25062: log10_cal = 16'b0000010110001110;
            15'd25063: log10_cal = 16'b0000010110001110;
            15'd25064: log10_cal = 16'b0000010110001110;
            15'd25065: log10_cal = 16'b0000010110001110;
            15'd25066: log10_cal = 16'b0000010110001110;
            15'd25067: log10_cal = 16'b0000010110001110;
            15'd25068: log10_cal = 16'b0000010110001110;
            15'd25069: log10_cal = 16'b0000010110001110;
            15'd25070: log10_cal = 16'b0000010110001110;
            15'd25071: log10_cal = 16'b0000010110001110;
            15'd25072: log10_cal = 16'b0000010110001110;
            15'd25073: log10_cal = 16'b0000010110001110;
            15'd25074: log10_cal = 16'b0000010110001110;
            15'd25075: log10_cal = 16'b0000010110001110;
            15'd25076: log10_cal = 16'b0000010110001110;
            15'd25077: log10_cal = 16'b0000010110001110;
            15'd25078: log10_cal = 16'b0000010110001110;
            15'd25079: log10_cal = 16'b0000010110001110;
            15'd25080: log10_cal = 16'b0000010110001110;
            15'd25081: log10_cal = 16'b0000010110001110;
            15'd25082: log10_cal = 16'b0000010110001110;
            15'd25083: log10_cal = 16'b0000010110001110;
            15'd25084: log10_cal = 16'b0000010110001110;
            15'd25085: log10_cal = 16'b0000010110001110;
            15'd25086: log10_cal = 16'b0000010110001110;
            15'd25087: log10_cal = 16'b0000010110001110;
            15'd25088: log10_cal = 16'b0000010110001110;
            15'd25089: log10_cal = 16'b0000010110001110;
            15'd25090: log10_cal = 16'b0000010110001110;
            15'd25091: log10_cal = 16'b0000010110001110;
            15'd25092: log10_cal = 16'b0000010110001110;
            15'd25093: log10_cal = 16'b0000010110001110;
            15'd25094: log10_cal = 16'b0000010110001110;
            15'd25095: log10_cal = 16'b0000010110001110;
            15'd25096: log10_cal = 16'b0000010110001110;
            15'd25097: log10_cal = 16'b0000010110001110;
            15'd25098: log10_cal = 16'b0000010110001110;
            15'd25099: log10_cal = 16'b0000010110001110;
            15'd25100: log10_cal = 16'b0000010110001110;
            15'd25101: log10_cal = 16'b0000010110001110;
            15'd25102: log10_cal = 16'b0000010110001110;
            15'd25103: log10_cal = 16'b0000010110001110;
            15'd25104: log10_cal = 16'b0000010110001110;
            15'd25105: log10_cal = 16'b0000010110001110;
            15'd25106: log10_cal = 16'b0000010110001110;
            15'd25107: log10_cal = 16'b0000010110001110;
            15'd25108: log10_cal = 16'b0000010110001110;
            15'd25109: log10_cal = 16'b0000010110001110;
            15'd25110: log10_cal = 16'b0000010110001110;
            15'd25111: log10_cal = 16'b0000010110001110;
            15'd25112: log10_cal = 16'b0000010110001110;
            15'd25113: log10_cal = 16'b0000010110001110;
            15'd25114: log10_cal = 16'b0000010110001110;
            15'd25115: log10_cal = 16'b0000010110001110;
            15'd25116: log10_cal = 16'b0000010110001111;
            15'd25117: log10_cal = 16'b0000010110001111;
            15'd25118: log10_cal = 16'b0000010110001111;
            15'd25119: log10_cal = 16'b0000010110001111;
            15'd25120: log10_cal = 16'b0000010110001111;
            15'd25121: log10_cal = 16'b0000010110001111;
            15'd25122: log10_cal = 16'b0000010110001111;
            15'd25123: log10_cal = 16'b0000010110001111;
            15'd25124: log10_cal = 16'b0000010110001111;
            15'd25125: log10_cal = 16'b0000010110001111;
            15'd25126: log10_cal = 16'b0000010110001111;
            15'd25127: log10_cal = 16'b0000010110001111;
            15'd25128: log10_cal = 16'b0000010110001111;
            15'd25129: log10_cal = 16'b0000010110001111;
            15'd25130: log10_cal = 16'b0000010110001111;
            15'd25131: log10_cal = 16'b0000010110001111;
            15'd25132: log10_cal = 16'b0000010110001111;
            15'd25133: log10_cal = 16'b0000010110001111;
            15'd25134: log10_cal = 16'b0000010110001111;
            15'd25135: log10_cal = 16'b0000010110001111;
            15'd25136: log10_cal = 16'b0000010110001111;
            15'd25137: log10_cal = 16'b0000010110001111;
            15'd25138: log10_cal = 16'b0000010110001111;
            15'd25139: log10_cal = 16'b0000010110001111;
            15'd25140: log10_cal = 16'b0000010110001111;
            15'd25141: log10_cal = 16'b0000010110001111;
            15'd25142: log10_cal = 16'b0000010110001111;
            15'd25143: log10_cal = 16'b0000010110001111;
            15'd25144: log10_cal = 16'b0000010110001111;
            15'd25145: log10_cal = 16'b0000010110001111;
            15'd25146: log10_cal = 16'b0000010110001111;
            15'd25147: log10_cal = 16'b0000010110001111;
            15'd25148: log10_cal = 16'b0000010110001111;
            15'd25149: log10_cal = 16'b0000010110001111;
            15'd25150: log10_cal = 16'b0000010110001111;
            15'd25151: log10_cal = 16'b0000010110001111;
            15'd25152: log10_cal = 16'b0000010110001111;
            15'd25153: log10_cal = 16'b0000010110001111;
            15'd25154: log10_cal = 16'b0000010110001111;
            15'd25155: log10_cal = 16'b0000010110001111;
            15'd25156: log10_cal = 16'b0000010110001111;
            15'd25157: log10_cal = 16'b0000010110001111;
            15'd25158: log10_cal = 16'b0000010110001111;
            15'd25159: log10_cal = 16'b0000010110001111;
            15'd25160: log10_cal = 16'b0000010110001111;
            15'd25161: log10_cal = 16'b0000010110001111;
            15'd25162: log10_cal = 16'b0000010110001111;
            15'd25163: log10_cal = 16'b0000010110001111;
            15'd25164: log10_cal = 16'b0000010110001111;
            15'd25165: log10_cal = 16'b0000010110001111;
            15'd25166: log10_cal = 16'b0000010110001111;
            15'd25167: log10_cal = 16'b0000010110001111;
            15'd25168: log10_cal = 16'b0000010110001111;
            15'd25169: log10_cal = 16'b0000010110001111;
            15'd25170: log10_cal = 16'b0000010110001111;
            15'd25171: log10_cal = 16'b0000010110001111;
            15'd25172: log10_cal = 16'b0000010110001111;
            15'd25173: log10_cal = 16'b0000010110010000;
            15'd25174: log10_cal = 16'b0000010110010000;
            15'd25175: log10_cal = 16'b0000010110010000;
            15'd25176: log10_cal = 16'b0000010110010000;
            15'd25177: log10_cal = 16'b0000010110010000;
            15'd25178: log10_cal = 16'b0000010110010000;
            15'd25179: log10_cal = 16'b0000010110010000;
            15'd25180: log10_cal = 16'b0000010110010000;
            15'd25181: log10_cal = 16'b0000010110010000;
            15'd25182: log10_cal = 16'b0000010110010000;
            15'd25183: log10_cal = 16'b0000010110010000;
            15'd25184: log10_cal = 16'b0000010110010000;
            15'd25185: log10_cal = 16'b0000010110010000;
            15'd25186: log10_cal = 16'b0000010110010000;
            15'd25187: log10_cal = 16'b0000010110010000;
            15'd25188: log10_cal = 16'b0000010110010000;
            15'd25189: log10_cal = 16'b0000010110010000;
            15'd25190: log10_cal = 16'b0000010110010000;
            15'd25191: log10_cal = 16'b0000010110010000;
            15'd25192: log10_cal = 16'b0000010110010000;
            15'd25193: log10_cal = 16'b0000010110010000;
            15'd25194: log10_cal = 16'b0000010110010000;
            15'd25195: log10_cal = 16'b0000010110010000;
            15'd25196: log10_cal = 16'b0000010110010000;
            15'd25197: log10_cal = 16'b0000010110010000;
            15'd25198: log10_cal = 16'b0000010110010000;
            15'd25199: log10_cal = 16'b0000010110010000;
            15'd25200: log10_cal = 16'b0000010110010000;
            15'd25201: log10_cal = 16'b0000010110010000;
            15'd25202: log10_cal = 16'b0000010110010000;
            15'd25203: log10_cal = 16'b0000010110010000;
            15'd25204: log10_cal = 16'b0000010110010000;
            15'd25205: log10_cal = 16'b0000010110010000;
            15'd25206: log10_cal = 16'b0000010110010000;
            15'd25207: log10_cal = 16'b0000010110010000;
            15'd25208: log10_cal = 16'b0000010110010000;
            15'd25209: log10_cal = 16'b0000010110010000;
            15'd25210: log10_cal = 16'b0000010110010000;
            15'd25211: log10_cal = 16'b0000010110010000;
            15'd25212: log10_cal = 16'b0000010110010000;
            15'd25213: log10_cal = 16'b0000010110010000;
            15'd25214: log10_cal = 16'b0000010110010000;
            15'd25215: log10_cal = 16'b0000010110010000;
            15'd25216: log10_cal = 16'b0000010110010000;
            15'd25217: log10_cal = 16'b0000010110010000;
            15'd25218: log10_cal = 16'b0000010110010000;
            15'd25219: log10_cal = 16'b0000010110010000;
            15'd25220: log10_cal = 16'b0000010110010000;
            15'd25221: log10_cal = 16'b0000010110010000;
            15'd25222: log10_cal = 16'b0000010110010000;
            15'd25223: log10_cal = 16'b0000010110010000;
            15'd25224: log10_cal = 16'b0000010110010000;
            15'd25225: log10_cal = 16'b0000010110010000;
            15'd25226: log10_cal = 16'b0000010110010000;
            15'd25227: log10_cal = 16'b0000010110010000;
            15'd25228: log10_cal = 16'b0000010110010000;
            15'd25229: log10_cal = 16'b0000010110010000;
            15'd25230: log10_cal = 16'b0000010110010001;
            15'd25231: log10_cal = 16'b0000010110010001;
            15'd25232: log10_cal = 16'b0000010110010001;
            15'd25233: log10_cal = 16'b0000010110010001;
            15'd25234: log10_cal = 16'b0000010110010001;
            15'd25235: log10_cal = 16'b0000010110010001;
            15'd25236: log10_cal = 16'b0000010110010001;
            15'd25237: log10_cal = 16'b0000010110010001;
            15'd25238: log10_cal = 16'b0000010110010001;
            15'd25239: log10_cal = 16'b0000010110010001;
            15'd25240: log10_cal = 16'b0000010110010001;
            15'd25241: log10_cal = 16'b0000010110010001;
            15'd25242: log10_cal = 16'b0000010110010001;
            15'd25243: log10_cal = 16'b0000010110010001;
            15'd25244: log10_cal = 16'b0000010110010001;
            15'd25245: log10_cal = 16'b0000010110010001;
            15'd25246: log10_cal = 16'b0000010110010001;
            15'd25247: log10_cal = 16'b0000010110010001;
            15'd25248: log10_cal = 16'b0000010110010001;
            15'd25249: log10_cal = 16'b0000010110010001;
            15'd25250: log10_cal = 16'b0000010110010001;
            15'd25251: log10_cal = 16'b0000010110010001;
            15'd25252: log10_cal = 16'b0000010110010001;
            15'd25253: log10_cal = 16'b0000010110010001;
            15'd25254: log10_cal = 16'b0000010110010001;
            15'd25255: log10_cal = 16'b0000010110010001;
            15'd25256: log10_cal = 16'b0000010110010001;
            15'd25257: log10_cal = 16'b0000010110010001;
            15'd25258: log10_cal = 16'b0000010110010001;
            15'd25259: log10_cal = 16'b0000010110010001;
            15'd25260: log10_cal = 16'b0000010110010001;
            15'd25261: log10_cal = 16'b0000010110010001;
            15'd25262: log10_cal = 16'b0000010110010001;
            15'd25263: log10_cal = 16'b0000010110010001;
            15'd25264: log10_cal = 16'b0000010110010001;
            15'd25265: log10_cal = 16'b0000010110010001;
            15'd25266: log10_cal = 16'b0000010110010001;
            15'd25267: log10_cal = 16'b0000010110010001;
            15'd25268: log10_cal = 16'b0000010110010001;
            15'd25269: log10_cal = 16'b0000010110010001;
            15'd25270: log10_cal = 16'b0000010110010001;
            15'd25271: log10_cal = 16'b0000010110010001;
            15'd25272: log10_cal = 16'b0000010110010001;
            15'd25273: log10_cal = 16'b0000010110010001;
            15'd25274: log10_cal = 16'b0000010110010001;
            15'd25275: log10_cal = 16'b0000010110010001;
            15'd25276: log10_cal = 16'b0000010110010001;
            15'd25277: log10_cal = 16'b0000010110010001;
            15'd25278: log10_cal = 16'b0000010110010001;
            15'd25279: log10_cal = 16'b0000010110010001;
            15'd25280: log10_cal = 16'b0000010110010001;
            15'd25281: log10_cal = 16'b0000010110010001;
            15'd25282: log10_cal = 16'b0000010110010001;
            15'd25283: log10_cal = 16'b0000010110010001;
            15'd25284: log10_cal = 16'b0000010110010001;
            15'd25285: log10_cal = 16'b0000010110010001;
            15'd25286: log10_cal = 16'b0000010110010010;
            15'd25287: log10_cal = 16'b0000010110010010;
            15'd25288: log10_cal = 16'b0000010110010010;
            15'd25289: log10_cal = 16'b0000010110010010;
            15'd25290: log10_cal = 16'b0000010110010010;
            15'd25291: log10_cal = 16'b0000010110010010;
            15'd25292: log10_cal = 16'b0000010110010010;
            15'd25293: log10_cal = 16'b0000010110010010;
            15'd25294: log10_cal = 16'b0000010110010010;
            15'd25295: log10_cal = 16'b0000010110010010;
            15'd25296: log10_cal = 16'b0000010110010010;
            15'd25297: log10_cal = 16'b0000010110010010;
            15'd25298: log10_cal = 16'b0000010110010010;
            15'd25299: log10_cal = 16'b0000010110010010;
            15'd25300: log10_cal = 16'b0000010110010010;
            15'd25301: log10_cal = 16'b0000010110010010;
            15'd25302: log10_cal = 16'b0000010110010010;
            15'd25303: log10_cal = 16'b0000010110010010;
            15'd25304: log10_cal = 16'b0000010110010010;
            15'd25305: log10_cal = 16'b0000010110010010;
            15'd25306: log10_cal = 16'b0000010110010010;
            15'd25307: log10_cal = 16'b0000010110010010;
            15'd25308: log10_cal = 16'b0000010110010010;
            15'd25309: log10_cal = 16'b0000010110010010;
            15'd25310: log10_cal = 16'b0000010110010010;
            15'd25311: log10_cal = 16'b0000010110010010;
            15'd25312: log10_cal = 16'b0000010110010010;
            15'd25313: log10_cal = 16'b0000010110010010;
            15'd25314: log10_cal = 16'b0000010110010010;
            15'd25315: log10_cal = 16'b0000010110010010;
            15'd25316: log10_cal = 16'b0000010110010010;
            15'd25317: log10_cal = 16'b0000010110010010;
            15'd25318: log10_cal = 16'b0000010110010010;
            15'd25319: log10_cal = 16'b0000010110010010;
            15'd25320: log10_cal = 16'b0000010110010010;
            15'd25321: log10_cal = 16'b0000010110010010;
            15'd25322: log10_cal = 16'b0000010110010010;
            15'd25323: log10_cal = 16'b0000010110010010;
            15'd25324: log10_cal = 16'b0000010110010010;
            15'd25325: log10_cal = 16'b0000010110010010;
            15'd25326: log10_cal = 16'b0000010110010010;
            15'd25327: log10_cal = 16'b0000010110010010;
            15'd25328: log10_cal = 16'b0000010110010010;
            15'd25329: log10_cal = 16'b0000010110010010;
            15'd25330: log10_cal = 16'b0000010110010010;
            15'd25331: log10_cal = 16'b0000010110010010;
            15'd25332: log10_cal = 16'b0000010110010010;
            15'd25333: log10_cal = 16'b0000010110010010;
            15'd25334: log10_cal = 16'b0000010110010010;
            15'd25335: log10_cal = 16'b0000010110010010;
            15'd25336: log10_cal = 16'b0000010110010010;
            15'd25337: log10_cal = 16'b0000010110010010;
            15'd25338: log10_cal = 16'b0000010110010010;
            15'd25339: log10_cal = 16'b0000010110010010;
            15'd25340: log10_cal = 16'b0000010110010010;
            15'd25341: log10_cal = 16'b0000010110010010;
            15'd25342: log10_cal = 16'b0000010110010010;
            15'd25343: log10_cal = 16'b0000010110010011;
            15'd25344: log10_cal = 16'b0000010110010011;
            15'd25345: log10_cal = 16'b0000010110010011;
            15'd25346: log10_cal = 16'b0000010110010011;
            15'd25347: log10_cal = 16'b0000010110010011;
            15'd25348: log10_cal = 16'b0000010110010011;
            15'd25349: log10_cal = 16'b0000010110010011;
            15'd25350: log10_cal = 16'b0000010110010011;
            15'd25351: log10_cal = 16'b0000010110010011;
            15'd25352: log10_cal = 16'b0000010110010011;
            15'd25353: log10_cal = 16'b0000010110010011;
            15'd25354: log10_cal = 16'b0000010110010011;
            15'd25355: log10_cal = 16'b0000010110010011;
            15'd25356: log10_cal = 16'b0000010110010011;
            15'd25357: log10_cal = 16'b0000010110010011;
            15'd25358: log10_cal = 16'b0000010110010011;
            15'd25359: log10_cal = 16'b0000010110010011;
            15'd25360: log10_cal = 16'b0000010110010011;
            15'd25361: log10_cal = 16'b0000010110010011;
            15'd25362: log10_cal = 16'b0000010110010011;
            15'd25363: log10_cal = 16'b0000010110010011;
            15'd25364: log10_cal = 16'b0000010110010011;
            15'd25365: log10_cal = 16'b0000010110010011;
            15'd25366: log10_cal = 16'b0000010110010011;
            15'd25367: log10_cal = 16'b0000010110010011;
            15'd25368: log10_cal = 16'b0000010110010011;
            15'd25369: log10_cal = 16'b0000010110010011;
            15'd25370: log10_cal = 16'b0000010110010011;
            15'd25371: log10_cal = 16'b0000010110010011;
            15'd25372: log10_cal = 16'b0000010110010011;
            15'd25373: log10_cal = 16'b0000010110010011;
            15'd25374: log10_cal = 16'b0000010110010011;
            15'd25375: log10_cal = 16'b0000010110010011;
            15'd25376: log10_cal = 16'b0000010110010011;
            15'd25377: log10_cal = 16'b0000010110010011;
            15'd25378: log10_cal = 16'b0000010110010011;
            15'd25379: log10_cal = 16'b0000010110010011;
            15'd25380: log10_cal = 16'b0000010110010011;
            15'd25381: log10_cal = 16'b0000010110010011;
            15'd25382: log10_cal = 16'b0000010110010011;
            15'd25383: log10_cal = 16'b0000010110010011;
            15'd25384: log10_cal = 16'b0000010110010011;
            15'd25385: log10_cal = 16'b0000010110010011;
            15'd25386: log10_cal = 16'b0000010110010011;
            15'd25387: log10_cal = 16'b0000010110010011;
            15'd25388: log10_cal = 16'b0000010110010011;
            15'd25389: log10_cal = 16'b0000010110010011;
            15'd25390: log10_cal = 16'b0000010110010011;
            15'd25391: log10_cal = 16'b0000010110010011;
            15'd25392: log10_cal = 16'b0000010110010011;
            15'd25393: log10_cal = 16'b0000010110010011;
            15'd25394: log10_cal = 16'b0000010110010011;
            15'd25395: log10_cal = 16'b0000010110010011;
            15'd25396: log10_cal = 16'b0000010110010011;
            15'd25397: log10_cal = 16'b0000010110010011;
            15'd25398: log10_cal = 16'b0000010110010011;
            15'd25399: log10_cal = 16'b0000010110010011;
            15'd25400: log10_cal = 16'b0000010110010100;
            15'd25401: log10_cal = 16'b0000010110010100;
            15'd25402: log10_cal = 16'b0000010110010100;
            15'd25403: log10_cal = 16'b0000010110010100;
            15'd25404: log10_cal = 16'b0000010110010100;
            15'd25405: log10_cal = 16'b0000010110010100;
            15'd25406: log10_cal = 16'b0000010110010100;
            15'd25407: log10_cal = 16'b0000010110010100;
            15'd25408: log10_cal = 16'b0000010110010100;
            15'd25409: log10_cal = 16'b0000010110010100;
            15'd25410: log10_cal = 16'b0000010110010100;
            15'd25411: log10_cal = 16'b0000010110010100;
            15'd25412: log10_cal = 16'b0000010110010100;
            15'd25413: log10_cal = 16'b0000010110010100;
            15'd25414: log10_cal = 16'b0000010110010100;
            15'd25415: log10_cal = 16'b0000010110010100;
            15'd25416: log10_cal = 16'b0000010110010100;
            15'd25417: log10_cal = 16'b0000010110010100;
            15'd25418: log10_cal = 16'b0000010110010100;
            15'd25419: log10_cal = 16'b0000010110010100;
            15'd25420: log10_cal = 16'b0000010110010100;
            15'd25421: log10_cal = 16'b0000010110010100;
            15'd25422: log10_cal = 16'b0000010110010100;
            15'd25423: log10_cal = 16'b0000010110010100;
            15'd25424: log10_cal = 16'b0000010110010100;
            15'd25425: log10_cal = 16'b0000010110010100;
            15'd25426: log10_cal = 16'b0000010110010100;
            15'd25427: log10_cal = 16'b0000010110010100;
            15'd25428: log10_cal = 16'b0000010110010100;
            15'd25429: log10_cal = 16'b0000010110010100;
            15'd25430: log10_cal = 16'b0000010110010100;
            15'd25431: log10_cal = 16'b0000010110010100;
            15'd25432: log10_cal = 16'b0000010110010100;
            15'd25433: log10_cal = 16'b0000010110010100;
            15'd25434: log10_cal = 16'b0000010110010100;
            15'd25435: log10_cal = 16'b0000010110010100;
            15'd25436: log10_cal = 16'b0000010110010100;
            15'd25437: log10_cal = 16'b0000010110010100;
            15'd25438: log10_cal = 16'b0000010110010100;
            15'd25439: log10_cal = 16'b0000010110010100;
            15'd25440: log10_cal = 16'b0000010110010100;
            15'd25441: log10_cal = 16'b0000010110010100;
            15'd25442: log10_cal = 16'b0000010110010100;
            15'd25443: log10_cal = 16'b0000010110010100;
            15'd25444: log10_cal = 16'b0000010110010100;
            15'd25445: log10_cal = 16'b0000010110010100;
            15'd25446: log10_cal = 16'b0000010110010100;
            15'd25447: log10_cal = 16'b0000010110010100;
            15'd25448: log10_cal = 16'b0000010110010100;
            15'd25449: log10_cal = 16'b0000010110010100;
            15'd25450: log10_cal = 16'b0000010110010100;
            15'd25451: log10_cal = 16'b0000010110010100;
            15'd25452: log10_cal = 16'b0000010110010100;
            15'd25453: log10_cal = 16'b0000010110010100;
            15'd25454: log10_cal = 16'b0000010110010100;
            15'd25455: log10_cal = 16'b0000010110010100;
            15'd25456: log10_cal = 16'b0000010110010100;
            15'd25457: log10_cal = 16'b0000010110010100;
            15'd25458: log10_cal = 16'b0000010110010101;
            15'd25459: log10_cal = 16'b0000010110010101;
            15'd25460: log10_cal = 16'b0000010110010101;
            15'd25461: log10_cal = 16'b0000010110010101;
            15'd25462: log10_cal = 16'b0000010110010101;
            15'd25463: log10_cal = 16'b0000010110010101;
            15'd25464: log10_cal = 16'b0000010110010101;
            15'd25465: log10_cal = 16'b0000010110010101;
            15'd25466: log10_cal = 16'b0000010110010101;
            15'd25467: log10_cal = 16'b0000010110010101;
            15'd25468: log10_cal = 16'b0000010110010101;
            15'd25469: log10_cal = 16'b0000010110010101;
            15'd25470: log10_cal = 16'b0000010110010101;
            15'd25471: log10_cal = 16'b0000010110010101;
            15'd25472: log10_cal = 16'b0000010110010101;
            15'd25473: log10_cal = 16'b0000010110010101;
            15'd25474: log10_cal = 16'b0000010110010101;
            15'd25475: log10_cal = 16'b0000010110010101;
            15'd25476: log10_cal = 16'b0000010110010101;
            15'd25477: log10_cal = 16'b0000010110010101;
            15'd25478: log10_cal = 16'b0000010110010101;
            15'd25479: log10_cal = 16'b0000010110010101;
            15'd25480: log10_cal = 16'b0000010110010101;
            15'd25481: log10_cal = 16'b0000010110010101;
            15'd25482: log10_cal = 16'b0000010110010101;
            15'd25483: log10_cal = 16'b0000010110010101;
            15'd25484: log10_cal = 16'b0000010110010101;
            15'd25485: log10_cal = 16'b0000010110010101;
            15'd25486: log10_cal = 16'b0000010110010101;
            15'd25487: log10_cal = 16'b0000010110010101;
            15'd25488: log10_cal = 16'b0000010110010101;
            15'd25489: log10_cal = 16'b0000010110010101;
            15'd25490: log10_cal = 16'b0000010110010101;
            15'd25491: log10_cal = 16'b0000010110010101;
            15'd25492: log10_cal = 16'b0000010110010101;
            15'd25493: log10_cal = 16'b0000010110010101;
            15'd25494: log10_cal = 16'b0000010110010101;
            15'd25495: log10_cal = 16'b0000010110010101;
            15'd25496: log10_cal = 16'b0000010110010101;
            15'd25497: log10_cal = 16'b0000010110010101;
            15'd25498: log10_cal = 16'b0000010110010101;
            15'd25499: log10_cal = 16'b0000010110010101;
            15'd25500: log10_cal = 16'b0000010110010101;
            15'd25501: log10_cal = 16'b0000010110010101;
            15'd25502: log10_cal = 16'b0000010110010101;
            15'd25503: log10_cal = 16'b0000010110010101;
            15'd25504: log10_cal = 16'b0000010110010101;
            15'd25505: log10_cal = 16'b0000010110010101;
            15'd25506: log10_cal = 16'b0000010110010101;
            15'd25507: log10_cal = 16'b0000010110010101;
            15'd25508: log10_cal = 16'b0000010110010101;
            15'd25509: log10_cal = 16'b0000010110010101;
            15'd25510: log10_cal = 16'b0000010110010101;
            15'd25511: log10_cal = 16'b0000010110010101;
            15'd25512: log10_cal = 16'b0000010110010101;
            15'd25513: log10_cal = 16'b0000010110010101;
            15'd25514: log10_cal = 16'b0000010110010101;
            15'd25515: log10_cal = 16'b0000010110010110;
            15'd25516: log10_cal = 16'b0000010110010110;
            15'd25517: log10_cal = 16'b0000010110010110;
            15'd25518: log10_cal = 16'b0000010110010110;
            15'd25519: log10_cal = 16'b0000010110010110;
            15'd25520: log10_cal = 16'b0000010110010110;
            15'd25521: log10_cal = 16'b0000010110010110;
            15'd25522: log10_cal = 16'b0000010110010110;
            15'd25523: log10_cal = 16'b0000010110010110;
            15'd25524: log10_cal = 16'b0000010110010110;
            15'd25525: log10_cal = 16'b0000010110010110;
            15'd25526: log10_cal = 16'b0000010110010110;
            15'd25527: log10_cal = 16'b0000010110010110;
            15'd25528: log10_cal = 16'b0000010110010110;
            15'd25529: log10_cal = 16'b0000010110010110;
            15'd25530: log10_cal = 16'b0000010110010110;
            15'd25531: log10_cal = 16'b0000010110010110;
            15'd25532: log10_cal = 16'b0000010110010110;
            15'd25533: log10_cal = 16'b0000010110010110;
            15'd25534: log10_cal = 16'b0000010110010110;
            15'd25535: log10_cal = 16'b0000010110010110;
            15'd25536: log10_cal = 16'b0000010110010110;
            15'd25537: log10_cal = 16'b0000010110010110;
            15'd25538: log10_cal = 16'b0000010110010110;
            15'd25539: log10_cal = 16'b0000010110010110;
            15'd25540: log10_cal = 16'b0000010110010110;
            15'd25541: log10_cal = 16'b0000010110010110;
            15'd25542: log10_cal = 16'b0000010110010110;
            15'd25543: log10_cal = 16'b0000010110010110;
            15'd25544: log10_cal = 16'b0000010110010110;
            15'd25545: log10_cal = 16'b0000010110010110;
            15'd25546: log10_cal = 16'b0000010110010110;
            15'd25547: log10_cal = 16'b0000010110010110;
            15'd25548: log10_cal = 16'b0000010110010110;
            15'd25549: log10_cal = 16'b0000010110010110;
            15'd25550: log10_cal = 16'b0000010110010110;
            15'd25551: log10_cal = 16'b0000010110010110;
            15'd25552: log10_cal = 16'b0000010110010110;
            15'd25553: log10_cal = 16'b0000010110010110;
            15'd25554: log10_cal = 16'b0000010110010110;
            15'd25555: log10_cal = 16'b0000010110010110;
            15'd25556: log10_cal = 16'b0000010110010110;
            15'd25557: log10_cal = 16'b0000010110010110;
            15'd25558: log10_cal = 16'b0000010110010110;
            15'd25559: log10_cal = 16'b0000010110010110;
            15'd25560: log10_cal = 16'b0000010110010110;
            15'd25561: log10_cal = 16'b0000010110010110;
            15'd25562: log10_cal = 16'b0000010110010110;
            15'd25563: log10_cal = 16'b0000010110010110;
            15'd25564: log10_cal = 16'b0000010110010110;
            15'd25565: log10_cal = 16'b0000010110010110;
            15'd25566: log10_cal = 16'b0000010110010110;
            15'd25567: log10_cal = 16'b0000010110010110;
            15'd25568: log10_cal = 16'b0000010110010110;
            15'd25569: log10_cal = 16'b0000010110010110;
            15'd25570: log10_cal = 16'b0000010110010110;
            15'd25571: log10_cal = 16'b0000010110010110;
            15'd25572: log10_cal = 16'b0000010110010111;
            15'd25573: log10_cal = 16'b0000010110010111;
            15'd25574: log10_cal = 16'b0000010110010111;
            15'd25575: log10_cal = 16'b0000010110010111;
            15'd25576: log10_cal = 16'b0000010110010111;
            15'd25577: log10_cal = 16'b0000010110010111;
            15'd25578: log10_cal = 16'b0000010110010111;
            15'd25579: log10_cal = 16'b0000010110010111;
            15'd25580: log10_cal = 16'b0000010110010111;
            15'd25581: log10_cal = 16'b0000010110010111;
            15'd25582: log10_cal = 16'b0000010110010111;
            15'd25583: log10_cal = 16'b0000010110010111;
            15'd25584: log10_cal = 16'b0000010110010111;
            15'd25585: log10_cal = 16'b0000010110010111;
            15'd25586: log10_cal = 16'b0000010110010111;
            15'd25587: log10_cal = 16'b0000010110010111;
            15'd25588: log10_cal = 16'b0000010110010111;
            15'd25589: log10_cal = 16'b0000010110010111;
            15'd25590: log10_cal = 16'b0000010110010111;
            15'd25591: log10_cal = 16'b0000010110010111;
            15'd25592: log10_cal = 16'b0000010110010111;
            15'd25593: log10_cal = 16'b0000010110010111;
            15'd25594: log10_cal = 16'b0000010110010111;
            15'd25595: log10_cal = 16'b0000010110010111;
            15'd25596: log10_cal = 16'b0000010110010111;
            15'd25597: log10_cal = 16'b0000010110010111;
            15'd25598: log10_cal = 16'b0000010110010111;
            15'd25599: log10_cal = 16'b0000010110010111;
            15'd25600: log10_cal = 16'b0000010110010111;
            15'd25601: log10_cal = 16'b0000010110010111;
            15'd25602: log10_cal = 16'b0000010110010111;
            15'd25603: log10_cal = 16'b0000010110010111;
            15'd25604: log10_cal = 16'b0000010110010111;
            15'd25605: log10_cal = 16'b0000010110010111;
            15'd25606: log10_cal = 16'b0000010110010111;
            15'd25607: log10_cal = 16'b0000010110010111;
            15'd25608: log10_cal = 16'b0000010110010111;
            15'd25609: log10_cal = 16'b0000010110010111;
            15'd25610: log10_cal = 16'b0000010110010111;
            15'd25611: log10_cal = 16'b0000010110010111;
            15'd25612: log10_cal = 16'b0000010110010111;
            15'd25613: log10_cal = 16'b0000010110010111;
            15'd25614: log10_cal = 16'b0000010110010111;
            15'd25615: log10_cal = 16'b0000010110010111;
            15'd25616: log10_cal = 16'b0000010110010111;
            15'd25617: log10_cal = 16'b0000010110010111;
            15'd25618: log10_cal = 16'b0000010110010111;
            15'd25619: log10_cal = 16'b0000010110010111;
            15'd25620: log10_cal = 16'b0000010110010111;
            15'd25621: log10_cal = 16'b0000010110010111;
            15'd25622: log10_cal = 16'b0000010110010111;
            15'd25623: log10_cal = 16'b0000010110010111;
            15'd25624: log10_cal = 16'b0000010110010111;
            15'd25625: log10_cal = 16'b0000010110010111;
            15'd25626: log10_cal = 16'b0000010110010111;
            15'd25627: log10_cal = 16'b0000010110010111;
            15'd25628: log10_cal = 16'b0000010110010111;
            15'd25629: log10_cal = 16'b0000010110010111;
            15'd25630: log10_cal = 16'b0000010110011000;
            15'd25631: log10_cal = 16'b0000010110011000;
            15'd25632: log10_cal = 16'b0000010110011000;
            15'd25633: log10_cal = 16'b0000010110011000;
            15'd25634: log10_cal = 16'b0000010110011000;
            15'd25635: log10_cal = 16'b0000010110011000;
            15'd25636: log10_cal = 16'b0000010110011000;
            15'd25637: log10_cal = 16'b0000010110011000;
            15'd25638: log10_cal = 16'b0000010110011000;
            15'd25639: log10_cal = 16'b0000010110011000;
            15'd25640: log10_cal = 16'b0000010110011000;
            15'd25641: log10_cal = 16'b0000010110011000;
            15'd25642: log10_cal = 16'b0000010110011000;
            15'd25643: log10_cal = 16'b0000010110011000;
            15'd25644: log10_cal = 16'b0000010110011000;
            15'd25645: log10_cal = 16'b0000010110011000;
            15'd25646: log10_cal = 16'b0000010110011000;
            15'd25647: log10_cal = 16'b0000010110011000;
            15'd25648: log10_cal = 16'b0000010110011000;
            15'd25649: log10_cal = 16'b0000010110011000;
            15'd25650: log10_cal = 16'b0000010110011000;
            15'd25651: log10_cal = 16'b0000010110011000;
            15'd25652: log10_cal = 16'b0000010110011000;
            15'd25653: log10_cal = 16'b0000010110011000;
            15'd25654: log10_cal = 16'b0000010110011000;
            15'd25655: log10_cal = 16'b0000010110011000;
            15'd25656: log10_cal = 16'b0000010110011000;
            15'd25657: log10_cal = 16'b0000010110011000;
            15'd25658: log10_cal = 16'b0000010110011000;
            15'd25659: log10_cal = 16'b0000010110011000;
            15'd25660: log10_cal = 16'b0000010110011000;
            15'd25661: log10_cal = 16'b0000010110011000;
            15'd25662: log10_cal = 16'b0000010110011000;
            15'd25663: log10_cal = 16'b0000010110011000;
            15'd25664: log10_cal = 16'b0000010110011000;
            15'd25665: log10_cal = 16'b0000010110011000;
            15'd25666: log10_cal = 16'b0000010110011000;
            15'd25667: log10_cal = 16'b0000010110011000;
            15'd25668: log10_cal = 16'b0000010110011000;
            15'd25669: log10_cal = 16'b0000010110011000;
            15'd25670: log10_cal = 16'b0000010110011000;
            15'd25671: log10_cal = 16'b0000010110011000;
            15'd25672: log10_cal = 16'b0000010110011000;
            15'd25673: log10_cal = 16'b0000010110011000;
            15'd25674: log10_cal = 16'b0000010110011000;
            15'd25675: log10_cal = 16'b0000010110011000;
            15'd25676: log10_cal = 16'b0000010110011000;
            15'd25677: log10_cal = 16'b0000010110011000;
            15'd25678: log10_cal = 16'b0000010110011000;
            15'd25679: log10_cal = 16'b0000010110011000;
            15'd25680: log10_cal = 16'b0000010110011000;
            15'd25681: log10_cal = 16'b0000010110011000;
            15'd25682: log10_cal = 16'b0000010110011000;
            15'd25683: log10_cal = 16'b0000010110011000;
            15'd25684: log10_cal = 16'b0000010110011000;
            15'd25685: log10_cal = 16'b0000010110011000;
            15'd25686: log10_cal = 16'b0000010110011000;
            15'd25687: log10_cal = 16'b0000010110011000;
            15'd25688: log10_cal = 16'b0000010110011001;
            15'd25689: log10_cal = 16'b0000010110011001;
            15'd25690: log10_cal = 16'b0000010110011001;
            15'd25691: log10_cal = 16'b0000010110011001;
            15'd25692: log10_cal = 16'b0000010110011001;
            15'd25693: log10_cal = 16'b0000010110011001;
            15'd25694: log10_cal = 16'b0000010110011001;
            15'd25695: log10_cal = 16'b0000010110011001;
            15'd25696: log10_cal = 16'b0000010110011001;
            15'd25697: log10_cal = 16'b0000010110011001;
            15'd25698: log10_cal = 16'b0000010110011001;
            15'd25699: log10_cal = 16'b0000010110011001;
            15'd25700: log10_cal = 16'b0000010110011001;
            15'd25701: log10_cal = 16'b0000010110011001;
            15'd25702: log10_cal = 16'b0000010110011001;
            15'd25703: log10_cal = 16'b0000010110011001;
            15'd25704: log10_cal = 16'b0000010110011001;
            15'd25705: log10_cal = 16'b0000010110011001;
            15'd25706: log10_cal = 16'b0000010110011001;
            15'd25707: log10_cal = 16'b0000010110011001;
            15'd25708: log10_cal = 16'b0000010110011001;
            15'd25709: log10_cal = 16'b0000010110011001;
            15'd25710: log10_cal = 16'b0000010110011001;
            15'd25711: log10_cal = 16'b0000010110011001;
            15'd25712: log10_cal = 16'b0000010110011001;
            15'd25713: log10_cal = 16'b0000010110011001;
            15'd25714: log10_cal = 16'b0000010110011001;
            15'd25715: log10_cal = 16'b0000010110011001;
            15'd25716: log10_cal = 16'b0000010110011001;
            15'd25717: log10_cal = 16'b0000010110011001;
            15'd25718: log10_cal = 16'b0000010110011001;
            15'd25719: log10_cal = 16'b0000010110011001;
            15'd25720: log10_cal = 16'b0000010110011001;
            15'd25721: log10_cal = 16'b0000010110011001;
            15'd25722: log10_cal = 16'b0000010110011001;
            15'd25723: log10_cal = 16'b0000010110011001;
            15'd25724: log10_cal = 16'b0000010110011001;
            15'd25725: log10_cal = 16'b0000010110011001;
            15'd25726: log10_cal = 16'b0000010110011001;
            15'd25727: log10_cal = 16'b0000010110011001;
            15'd25728: log10_cal = 16'b0000010110011001;
            15'd25729: log10_cal = 16'b0000010110011001;
            15'd25730: log10_cal = 16'b0000010110011001;
            15'd25731: log10_cal = 16'b0000010110011001;
            15'd25732: log10_cal = 16'b0000010110011001;
            15'd25733: log10_cal = 16'b0000010110011001;
            15'd25734: log10_cal = 16'b0000010110011001;
            15'd25735: log10_cal = 16'b0000010110011001;
            15'd25736: log10_cal = 16'b0000010110011001;
            15'd25737: log10_cal = 16'b0000010110011001;
            15'd25738: log10_cal = 16'b0000010110011001;
            15'd25739: log10_cal = 16'b0000010110011001;
            15'd25740: log10_cal = 16'b0000010110011001;
            15'd25741: log10_cal = 16'b0000010110011001;
            15'd25742: log10_cal = 16'b0000010110011001;
            15'd25743: log10_cal = 16'b0000010110011001;
            15'd25744: log10_cal = 16'b0000010110011001;
            15'd25745: log10_cal = 16'b0000010110011010;
            15'd25746: log10_cal = 16'b0000010110011010;
            15'd25747: log10_cal = 16'b0000010110011010;
            15'd25748: log10_cal = 16'b0000010110011010;
            15'd25749: log10_cal = 16'b0000010110011010;
            15'd25750: log10_cal = 16'b0000010110011010;
            15'd25751: log10_cal = 16'b0000010110011010;
            15'd25752: log10_cal = 16'b0000010110011010;
            15'd25753: log10_cal = 16'b0000010110011010;
            15'd25754: log10_cal = 16'b0000010110011010;
            15'd25755: log10_cal = 16'b0000010110011010;
            15'd25756: log10_cal = 16'b0000010110011010;
            15'd25757: log10_cal = 16'b0000010110011010;
            15'd25758: log10_cal = 16'b0000010110011010;
            15'd25759: log10_cal = 16'b0000010110011010;
            15'd25760: log10_cal = 16'b0000010110011010;
            15'd25761: log10_cal = 16'b0000010110011010;
            15'd25762: log10_cal = 16'b0000010110011010;
            15'd25763: log10_cal = 16'b0000010110011010;
            15'd25764: log10_cal = 16'b0000010110011010;
            15'd25765: log10_cal = 16'b0000010110011010;
            15'd25766: log10_cal = 16'b0000010110011010;
            15'd25767: log10_cal = 16'b0000010110011010;
            15'd25768: log10_cal = 16'b0000010110011010;
            15'd25769: log10_cal = 16'b0000010110011010;
            15'd25770: log10_cal = 16'b0000010110011010;
            15'd25771: log10_cal = 16'b0000010110011010;
            15'd25772: log10_cal = 16'b0000010110011010;
            15'd25773: log10_cal = 16'b0000010110011010;
            15'd25774: log10_cal = 16'b0000010110011010;
            15'd25775: log10_cal = 16'b0000010110011010;
            15'd25776: log10_cal = 16'b0000010110011010;
            15'd25777: log10_cal = 16'b0000010110011010;
            15'd25778: log10_cal = 16'b0000010110011010;
            15'd25779: log10_cal = 16'b0000010110011010;
            15'd25780: log10_cal = 16'b0000010110011010;
            15'd25781: log10_cal = 16'b0000010110011010;
            15'd25782: log10_cal = 16'b0000010110011010;
            15'd25783: log10_cal = 16'b0000010110011010;
            15'd25784: log10_cal = 16'b0000010110011010;
            15'd25785: log10_cal = 16'b0000010110011010;
            15'd25786: log10_cal = 16'b0000010110011010;
            15'd25787: log10_cal = 16'b0000010110011010;
            15'd25788: log10_cal = 16'b0000010110011010;
            15'd25789: log10_cal = 16'b0000010110011010;
            15'd25790: log10_cal = 16'b0000010110011010;
            15'd25791: log10_cal = 16'b0000010110011010;
            15'd25792: log10_cal = 16'b0000010110011010;
            15'd25793: log10_cal = 16'b0000010110011010;
            15'd25794: log10_cal = 16'b0000010110011010;
            15'd25795: log10_cal = 16'b0000010110011010;
            15'd25796: log10_cal = 16'b0000010110011010;
            15'd25797: log10_cal = 16'b0000010110011010;
            15'd25798: log10_cal = 16'b0000010110011010;
            15'd25799: log10_cal = 16'b0000010110011010;
            15'd25800: log10_cal = 16'b0000010110011010;
            15'd25801: log10_cal = 16'b0000010110011010;
            15'd25802: log10_cal = 16'b0000010110011010;
            15'd25803: log10_cal = 16'b0000010110011011;
            15'd25804: log10_cal = 16'b0000010110011011;
            15'd25805: log10_cal = 16'b0000010110011011;
            15'd25806: log10_cal = 16'b0000010110011011;
            15'd25807: log10_cal = 16'b0000010110011011;
            15'd25808: log10_cal = 16'b0000010110011011;
            15'd25809: log10_cal = 16'b0000010110011011;
            15'd25810: log10_cal = 16'b0000010110011011;
            15'd25811: log10_cal = 16'b0000010110011011;
            15'd25812: log10_cal = 16'b0000010110011011;
            15'd25813: log10_cal = 16'b0000010110011011;
            15'd25814: log10_cal = 16'b0000010110011011;
            15'd25815: log10_cal = 16'b0000010110011011;
            15'd25816: log10_cal = 16'b0000010110011011;
            15'd25817: log10_cal = 16'b0000010110011011;
            15'd25818: log10_cal = 16'b0000010110011011;
            15'd25819: log10_cal = 16'b0000010110011011;
            15'd25820: log10_cal = 16'b0000010110011011;
            15'd25821: log10_cal = 16'b0000010110011011;
            15'd25822: log10_cal = 16'b0000010110011011;
            15'd25823: log10_cal = 16'b0000010110011011;
            15'd25824: log10_cal = 16'b0000010110011011;
            15'd25825: log10_cal = 16'b0000010110011011;
            15'd25826: log10_cal = 16'b0000010110011011;
            15'd25827: log10_cal = 16'b0000010110011011;
            15'd25828: log10_cal = 16'b0000010110011011;
            15'd25829: log10_cal = 16'b0000010110011011;
            15'd25830: log10_cal = 16'b0000010110011011;
            15'd25831: log10_cal = 16'b0000010110011011;
            15'd25832: log10_cal = 16'b0000010110011011;
            15'd25833: log10_cal = 16'b0000010110011011;
            15'd25834: log10_cal = 16'b0000010110011011;
            15'd25835: log10_cal = 16'b0000010110011011;
            15'd25836: log10_cal = 16'b0000010110011011;
            15'd25837: log10_cal = 16'b0000010110011011;
            15'd25838: log10_cal = 16'b0000010110011011;
            15'd25839: log10_cal = 16'b0000010110011011;
            15'd25840: log10_cal = 16'b0000010110011011;
            15'd25841: log10_cal = 16'b0000010110011011;
            15'd25842: log10_cal = 16'b0000010110011011;
            15'd25843: log10_cal = 16'b0000010110011011;
            15'd25844: log10_cal = 16'b0000010110011011;
            15'd25845: log10_cal = 16'b0000010110011011;
            15'd25846: log10_cal = 16'b0000010110011011;
            15'd25847: log10_cal = 16'b0000010110011011;
            15'd25848: log10_cal = 16'b0000010110011011;
            15'd25849: log10_cal = 16'b0000010110011011;
            15'd25850: log10_cal = 16'b0000010110011011;
            15'd25851: log10_cal = 16'b0000010110011011;
            15'd25852: log10_cal = 16'b0000010110011011;
            15'd25853: log10_cal = 16'b0000010110011011;
            15'd25854: log10_cal = 16'b0000010110011011;
            15'd25855: log10_cal = 16'b0000010110011011;
            15'd25856: log10_cal = 16'b0000010110011011;
            15'd25857: log10_cal = 16'b0000010110011011;
            15'd25858: log10_cal = 16'b0000010110011011;
            15'd25859: log10_cal = 16'b0000010110011011;
            15'd25860: log10_cal = 16'b0000010110011011;
            15'd25861: log10_cal = 16'b0000010110011100;
            15'd25862: log10_cal = 16'b0000010110011100;
            15'd25863: log10_cal = 16'b0000010110011100;
            15'd25864: log10_cal = 16'b0000010110011100;
            15'd25865: log10_cal = 16'b0000010110011100;
            15'd25866: log10_cal = 16'b0000010110011100;
            15'd25867: log10_cal = 16'b0000010110011100;
            15'd25868: log10_cal = 16'b0000010110011100;
            15'd25869: log10_cal = 16'b0000010110011100;
            15'd25870: log10_cal = 16'b0000010110011100;
            15'd25871: log10_cal = 16'b0000010110011100;
            15'd25872: log10_cal = 16'b0000010110011100;
            15'd25873: log10_cal = 16'b0000010110011100;
            15'd25874: log10_cal = 16'b0000010110011100;
            15'd25875: log10_cal = 16'b0000010110011100;
            15'd25876: log10_cal = 16'b0000010110011100;
            15'd25877: log10_cal = 16'b0000010110011100;
            15'd25878: log10_cal = 16'b0000010110011100;
            15'd25879: log10_cal = 16'b0000010110011100;
            15'd25880: log10_cal = 16'b0000010110011100;
            15'd25881: log10_cal = 16'b0000010110011100;
            15'd25882: log10_cal = 16'b0000010110011100;
            15'd25883: log10_cal = 16'b0000010110011100;
            15'd25884: log10_cal = 16'b0000010110011100;
            15'd25885: log10_cal = 16'b0000010110011100;
            15'd25886: log10_cal = 16'b0000010110011100;
            15'd25887: log10_cal = 16'b0000010110011100;
            15'd25888: log10_cal = 16'b0000010110011100;
            15'd25889: log10_cal = 16'b0000010110011100;
            15'd25890: log10_cal = 16'b0000010110011100;
            15'd25891: log10_cal = 16'b0000010110011100;
            15'd25892: log10_cal = 16'b0000010110011100;
            15'd25893: log10_cal = 16'b0000010110011100;
            15'd25894: log10_cal = 16'b0000010110011100;
            15'd25895: log10_cal = 16'b0000010110011100;
            15'd25896: log10_cal = 16'b0000010110011100;
            15'd25897: log10_cal = 16'b0000010110011100;
            15'd25898: log10_cal = 16'b0000010110011100;
            15'd25899: log10_cal = 16'b0000010110011100;
            15'd25900: log10_cal = 16'b0000010110011100;
            15'd25901: log10_cal = 16'b0000010110011100;
            15'd25902: log10_cal = 16'b0000010110011100;
            15'd25903: log10_cal = 16'b0000010110011100;
            15'd25904: log10_cal = 16'b0000010110011100;
            15'd25905: log10_cal = 16'b0000010110011100;
            15'd25906: log10_cal = 16'b0000010110011100;
            15'd25907: log10_cal = 16'b0000010110011100;
            15'd25908: log10_cal = 16'b0000010110011100;
            15'd25909: log10_cal = 16'b0000010110011100;
            15'd25910: log10_cal = 16'b0000010110011100;
            15'd25911: log10_cal = 16'b0000010110011100;
            15'd25912: log10_cal = 16'b0000010110011100;
            15'd25913: log10_cal = 16'b0000010110011100;
            15'd25914: log10_cal = 16'b0000010110011100;
            15'd25915: log10_cal = 16'b0000010110011100;
            15'd25916: log10_cal = 16'b0000010110011100;
            15'd25917: log10_cal = 16'b0000010110011100;
            15'd25918: log10_cal = 16'b0000010110011100;
            15'd25919: log10_cal = 16'b0000010110011100;
            15'd25920: log10_cal = 16'b0000010110011101;
            15'd25921: log10_cal = 16'b0000010110011101;
            15'd25922: log10_cal = 16'b0000010110011101;
            15'd25923: log10_cal = 16'b0000010110011101;
            15'd25924: log10_cal = 16'b0000010110011101;
            15'd25925: log10_cal = 16'b0000010110011101;
            15'd25926: log10_cal = 16'b0000010110011101;
            15'd25927: log10_cal = 16'b0000010110011101;
            15'd25928: log10_cal = 16'b0000010110011101;
            15'd25929: log10_cal = 16'b0000010110011101;
            15'd25930: log10_cal = 16'b0000010110011101;
            15'd25931: log10_cal = 16'b0000010110011101;
            15'd25932: log10_cal = 16'b0000010110011101;
            15'd25933: log10_cal = 16'b0000010110011101;
            15'd25934: log10_cal = 16'b0000010110011101;
            15'd25935: log10_cal = 16'b0000010110011101;
            15'd25936: log10_cal = 16'b0000010110011101;
            15'd25937: log10_cal = 16'b0000010110011101;
            15'd25938: log10_cal = 16'b0000010110011101;
            15'd25939: log10_cal = 16'b0000010110011101;
            15'd25940: log10_cal = 16'b0000010110011101;
            15'd25941: log10_cal = 16'b0000010110011101;
            15'd25942: log10_cal = 16'b0000010110011101;
            15'd25943: log10_cal = 16'b0000010110011101;
            15'd25944: log10_cal = 16'b0000010110011101;
            15'd25945: log10_cal = 16'b0000010110011101;
            15'd25946: log10_cal = 16'b0000010110011101;
            15'd25947: log10_cal = 16'b0000010110011101;
            15'd25948: log10_cal = 16'b0000010110011101;
            15'd25949: log10_cal = 16'b0000010110011101;
            15'd25950: log10_cal = 16'b0000010110011101;
            15'd25951: log10_cal = 16'b0000010110011101;
            15'd25952: log10_cal = 16'b0000010110011101;
            15'd25953: log10_cal = 16'b0000010110011101;
            15'd25954: log10_cal = 16'b0000010110011101;
            15'd25955: log10_cal = 16'b0000010110011101;
            15'd25956: log10_cal = 16'b0000010110011101;
            15'd25957: log10_cal = 16'b0000010110011101;
            15'd25958: log10_cal = 16'b0000010110011101;
            15'd25959: log10_cal = 16'b0000010110011101;
            15'd25960: log10_cal = 16'b0000010110011101;
            15'd25961: log10_cal = 16'b0000010110011101;
            15'd25962: log10_cal = 16'b0000010110011101;
            15'd25963: log10_cal = 16'b0000010110011101;
            15'd25964: log10_cal = 16'b0000010110011101;
            15'd25965: log10_cal = 16'b0000010110011101;
            15'd25966: log10_cal = 16'b0000010110011101;
            15'd25967: log10_cal = 16'b0000010110011101;
            15'd25968: log10_cal = 16'b0000010110011101;
            15'd25969: log10_cal = 16'b0000010110011101;
            15'd25970: log10_cal = 16'b0000010110011101;
            15'd25971: log10_cal = 16'b0000010110011101;
            15'd25972: log10_cal = 16'b0000010110011101;
            15'd25973: log10_cal = 16'b0000010110011101;
            15'd25974: log10_cal = 16'b0000010110011101;
            15'd25975: log10_cal = 16'b0000010110011101;
            15'd25976: log10_cal = 16'b0000010110011101;
            15'd25977: log10_cal = 16'b0000010110011101;
            15'd25978: log10_cal = 16'b0000010110011110;
            15'd25979: log10_cal = 16'b0000010110011110;
            15'd25980: log10_cal = 16'b0000010110011110;
            15'd25981: log10_cal = 16'b0000010110011110;
            15'd25982: log10_cal = 16'b0000010110011110;
            15'd25983: log10_cal = 16'b0000010110011110;
            15'd25984: log10_cal = 16'b0000010110011110;
            15'd25985: log10_cal = 16'b0000010110011110;
            15'd25986: log10_cal = 16'b0000010110011110;
            15'd25987: log10_cal = 16'b0000010110011110;
            15'd25988: log10_cal = 16'b0000010110011110;
            15'd25989: log10_cal = 16'b0000010110011110;
            15'd25990: log10_cal = 16'b0000010110011110;
            15'd25991: log10_cal = 16'b0000010110011110;
            15'd25992: log10_cal = 16'b0000010110011110;
            15'd25993: log10_cal = 16'b0000010110011110;
            15'd25994: log10_cal = 16'b0000010110011110;
            15'd25995: log10_cal = 16'b0000010110011110;
            15'd25996: log10_cal = 16'b0000010110011110;
            15'd25997: log10_cal = 16'b0000010110011110;
            15'd25998: log10_cal = 16'b0000010110011110;
            15'd25999: log10_cal = 16'b0000010110011110;
            15'd26000: log10_cal = 16'b0000010110011110;
            15'd26001: log10_cal = 16'b0000010110011110;
            15'd26002: log10_cal = 16'b0000010110011110;
            15'd26003: log10_cal = 16'b0000010110011110;
            15'd26004: log10_cal = 16'b0000010110011110;
            15'd26005: log10_cal = 16'b0000010110011110;
            15'd26006: log10_cal = 16'b0000010110011110;
            15'd26007: log10_cal = 16'b0000010110011110;
            15'd26008: log10_cal = 16'b0000010110011110;
            15'd26009: log10_cal = 16'b0000010110011110;
            15'd26010: log10_cal = 16'b0000010110011110;
            15'd26011: log10_cal = 16'b0000010110011110;
            15'd26012: log10_cal = 16'b0000010110011110;
            15'd26013: log10_cal = 16'b0000010110011110;
            15'd26014: log10_cal = 16'b0000010110011110;
            15'd26015: log10_cal = 16'b0000010110011110;
            15'd26016: log10_cal = 16'b0000010110011110;
            15'd26017: log10_cal = 16'b0000010110011110;
            15'd26018: log10_cal = 16'b0000010110011110;
            15'd26019: log10_cal = 16'b0000010110011110;
            15'd26020: log10_cal = 16'b0000010110011110;
            15'd26021: log10_cal = 16'b0000010110011110;
            15'd26022: log10_cal = 16'b0000010110011110;
            15'd26023: log10_cal = 16'b0000010110011110;
            15'd26024: log10_cal = 16'b0000010110011110;
            15'd26025: log10_cal = 16'b0000010110011110;
            15'd26026: log10_cal = 16'b0000010110011110;
            15'd26027: log10_cal = 16'b0000010110011110;
            15'd26028: log10_cal = 16'b0000010110011110;
            15'd26029: log10_cal = 16'b0000010110011110;
            15'd26030: log10_cal = 16'b0000010110011110;
            15'd26031: log10_cal = 16'b0000010110011110;
            15'd26032: log10_cal = 16'b0000010110011110;
            15'd26033: log10_cal = 16'b0000010110011110;
            15'd26034: log10_cal = 16'b0000010110011110;
            15'd26035: log10_cal = 16'b0000010110011110;
            15'd26036: log10_cal = 16'b0000010110011111;
            15'd26037: log10_cal = 16'b0000010110011111;
            15'd26038: log10_cal = 16'b0000010110011111;
            15'd26039: log10_cal = 16'b0000010110011111;
            15'd26040: log10_cal = 16'b0000010110011111;
            15'd26041: log10_cal = 16'b0000010110011111;
            15'd26042: log10_cal = 16'b0000010110011111;
            15'd26043: log10_cal = 16'b0000010110011111;
            15'd26044: log10_cal = 16'b0000010110011111;
            15'd26045: log10_cal = 16'b0000010110011111;
            15'd26046: log10_cal = 16'b0000010110011111;
            15'd26047: log10_cal = 16'b0000010110011111;
            15'd26048: log10_cal = 16'b0000010110011111;
            15'd26049: log10_cal = 16'b0000010110011111;
            15'd26050: log10_cal = 16'b0000010110011111;
            15'd26051: log10_cal = 16'b0000010110011111;
            15'd26052: log10_cal = 16'b0000010110011111;
            15'd26053: log10_cal = 16'b0000010110011111;
            15'd26054: log10_cal = 16'b0000010110011111;
            15'd26055: log10_cal = 16'b0000010110011111;
            15'd26056: log10_cal = 16'b0000010110011111;
            15'd26057: log10_cal = 16'b0000010110011111;
            15'd26058: log10_cal = 16'b0000010110011111;
            15'd26059: log10_cal = 16'b0000010110011111;
            15'd26060: log10_cal = 16'b0000010110011111;
            15'd26061: log10_cal = 16'b0000010110011111;
            15'd26062: log10_cal = 16'b0000010110011111;
            15'd26063: log10_cal = 16'b0000010110011111;
            15'd26064: log10_cal = 16'b0000010110011111;
            15'd26065: log10_cal = 16'b0000010110011111;
            15'd26066: log10_cal = 16'b0000010110011111;
            15'd26067: log10_cal = 16'b0000010110011111;
            15'd26068: log10_cal = 16'b0000010110011111;
            15'd26069: log10_cal = 16'b0000010110011111;
            15'd26070: log10_cal = 16'b0000010110011111;
            15'd26071: log10_cal = 16'b0000010110011111;
            15'd26072: log10_cal = 16'b0000010110011111;
            15'd26073: log10_cal = 16'b0000010110011111;
            15'd26074: log10_cal = 16'b0000010110011111;
            15'd26075: log10_cal = 16'b0000010110011111;
            15'd26076: log10_cal = 16'b0000010110011111;
            15'd26077: log10_cal = 16'b0000010110011111;
            15'd26078: log10_cal = 16'b0000010110011111;
            15'd26079: log10_cal = 16'b0000010110011111;
            15'd26080: log10_cal = 16'b0000010110011111;
            15'd26081: log10_cal = 16'b0000010110011111;
            15'd26082: log10_cal = 16'b0000010110011111;
            15'd26083: log10_cal = 16'b0000010110011111;
            15'd26084: log10_cal = 16'b0000010110011111;
            15'd26085: log10_cal = 16'b0000010110011111;
            15'd26086: log10_cal = 16'b0000010110011111;
            15'd26087: log10_cal = 16'b0000010110011111;
            15'd26088: log10_cal = 16'b0000010110011111;
            15'd26089: log10_cal = 16'b0000010110011111;
            15'd26090: log10_cal = 16'b0000010110011111;
            15'd26091: log10_cal = 16'b0000010110011111;
            15'd26092: log10_cal = 16'b0000010110011111;
            15'd26093: log10_cal = 16'b0000010110011111;
            15'd26094: log10_cal = 16'b0000010110011111;
            15'd26095: log10_cal = 16'b0000010110100000;
            15'd26096: log10_cal = 16'b0000010110100000;
            15'd26097: log10_cal = 16'b0000010110100000;
            15'd26098: log10_cal = 16'b0000010110100000;
            15'd26099: log10_cal = 16'b0000010110100000;
            15'd26100: log10_cal = 16'b0000010110100000;
            15'd26101: log10_cal = 16'b0000010110100000;
            15'd26102: log10_cal = 16'b0000010110100000;
            15'd26103: log10_cal = 16'b0000010110100000;
            15'd26104: log10_cal = 16'b0000010110100000;
            15'd26105: log10_cal = 16'b0000010110100000;
            15'd26106: log10_cal = 16'b0000010110100000;
            15'd26107: log10_cal = 16'b0000010110100000;
            15'd26108: log10_cal = 16'b0000010110100000;
            15'd26109: log10_cal = 16'b0000010110100000;
            15'd26110: log10_cal = 16'b0000010110100000;
            15'd26111: log10_cal = 16'b0000010110100000;
            15'd26112: log10_cal = 16'b0000010110100000;
            15'd26113: log10_cal = 16'b0000010110100000;
            15'd26114: log10_cal = 16'b0000010110100000;
            15'd26115: log10_cal = 16'b0000010110100000;
            15'd26116: log10_cal = 16'b0000010110100000;
            15'd26117: log10_cal = 16'b0000010110100000;
            15'd26118: log10_cal = 16'b0000010110100000;
            15'd26119: log10_cal = 16'b0000010110100000;
            15'd26120: log10_cal = 16'b0000010110100000;
            15'd26121: log10_cal = 16'b0000010110100000;
            15'd26122: log10_cal = 16'b0000010110100000;
            15'd26123: log10_cal = 16'b0000010110100000;
            15'd26124: log10_cal = 16'b0000010110100000;
            15'd26125: log10_cal = 16'b0000010110100000;
            15'd26126: log10_cal = 16'b0000010110100000;
            15'd26127: log10_cal = 16'b0000010110100000;
            15'd26128: log10_cal = 16'b0000010110100000;
            15'd26129: log10_cal = 16'b0000010110100000;
            15'd26130: log10_cal = 16'b0000010110100000;
            15'd26131: log10_cal = 16'b0000010110100000;
            15'd26132: log10_cal = 16'b0000010110100000;
            15'd26133: log10_cal = 16'b0000010110100000;
            15'd26134: log10_cal = 16'b0000010110100000;
            15'd26135: log10_cal = 16'b0000010110100000;
            15'd26136: log10_cal = 16'b0000010110100000;
            15'd26137: log10_cal = 16'b0000010110100000;
            15'd26138: log10_cal = 16'b0000010110100000;
            15'd26139: log10_cal = 16'b0000010110100000;
            15'd26140: log10_cal = 16'b0000010110100000;
            15'd26141: log10_cal = 16'b0000010110100000;
            15'd26142: log10_cal = 16'b0000010110100000;
            15'd26143: log10_cal = 16'b0000010110100000;
            15'd26144: log10_cal = 16'b0000010110100000;
            15'd26145: log10_cal = 16'b0000010110100000;
            15'd26146: log10_cal = 16'b0000010110100000;
            15'd26147: log10_cal = 16'b0000010110100000;
            15'd26148: log10_cal = 16'b0000010110100000;
            15'd26149: log10_cal = 16'b0000010110100000;
            15'd26150: log10_cal = 16'b0000010110100000;
            15'd26151: log10_cal = 16'b0000010110100000;
            15'd26152: log10_cal = 16'b0000010110100000;
            15'd26153: log10_cal = 16'b0000010110100000;
            15'd26154: log10_cal = 16'b0000010110100001;
            15'd26155: log10_cal = 16'b0000010110100001;
            15'd26156: log10_cal = 16'b0000010110100001;
            15'd26157: log10_cal = 16'b0000010110100001;
            15'd26158: log10_cal = 16'b0000010110100001;
            15'd26159: log10_cal = 16'b0000010110100001;
            15'd26160: log10_cal = 16'b0000010110100001;
            15'd26161: log10_cal = 16'b0000010110100001;
            15'd26162: log10_cal = 16'b0000010110100001;
            15'd26163: log10_cal = 16'b0000010110100001;
            15'd26164: log10_cal = 16'b0000010110100001;
            15'd26165: log10_cal = 16'b0000010110100001;
            15'd26166: log10_cal = 16'b0000010110100001;
            15'd26167: log10_cal = 16'b0000010110100001;
            15'd26168: log10_cal = 16'b0000010110100001;
            15'd26169: log10_cal = 16'b0000010110100001;
            15'd26170: log10_cal = 16'b0000010110100001;
            15'd26171: log10_cal = 16'b0000010110100001;
            15'd26172: log10_cal = 16'b0000010110100001;
            15'd26173: log10_cal = 16'b0000010110100001;
            15'd26174: log10_cal = 16'b0000010110100001;
            15'd26175: log10_cal = 16'b0000010110100001;
            15'd26176: log10_cal = 16'b0000010110100001;
            15'd26177: log10_cal = 16'b0000010110100001;
            15'd26178: log10_cal = 16'b0000010110100001;
            15'd26179: log10_cal = 16'b0000010110100001;
            15'd26180: log10_cal = 16'b0000010110100001;
            15'd26181: log10_cal = 16'b0000010110100001;
            15'd26182: log10_cal = 16'b0000010110100001;
            15'd26183: log10_cal = 16'b0000010110100001;
            15'd26184: log10_cal = 16'b0000010110100001;
            15'd26185: log10_cal = 16'b0000010110100001;
            15'd26186: log10_cal = 16'b0000010110100001;
            15'd26187: log10_cal = 16'b0000010110100001;
            15'd26188: log10_cal = 16'b0000010110100001;
            15'd26189: log10_cal = 16'b0000010110100001;
            15'd26190: log10_cal = 16'b0000010110100001;
            15'd26191: log10_cal = 16'b0000010110100001;
            15'd26192: log10_cal = 16'b0000010110100001;
            15'd26193: log10_cal = 16'b0000010110100001;
            15'd26194: log10_cal = 16'b0000010110100001;
            15'd26195: log10_cal = 16'b0000010110100001;
            15'd26196: log10_cal = 16'b0000010110100001;
            15'd26197: log10_cal = 16'b0000010110100001;
            15'd26198: log10_cal = 16'b0000010110100001;
            15'd26199: log10_cal = 16'b0000010110100001;
            15'd26200: log10_cal = 16'b0000010110100001;
            15'd26201: log10_cal = 16'b0000010110100001;
            15'd26202: log10_cal = 16'b0000010110100001;
            15'd26203: log10_cal = 16'b0000010110100001;
            15'd26204: log10_cal = 16'b0000010110100001;
            15'd26205: log10_cal = 16'b0000010110100001;
            15'd26206: log10_cal = 16'b0000010110100001;
            15'd26207: log10_cal = 16'b0000010110100001;
            15'd26208: log10_cal = 16'b0000010110100001;
            15'd26209: log10_cal = 16'b0000010110100001;
            15'd26210: log10_cal = 16'b0000010110100001;
            15'd26211: log10_cal = 16'b0000010110100001;
            15'd26212: log10_cal = 16'b0000010110100001;
            15'd26213: log10_cal = 16'b0000010110100010;
            15'd26214: log10_cal = 16'b0000010110100010;
            15'd26215: log10_cal = 16'b0000010110100010;
            15'd26216: log10_cal = 16'b0000010110100010;
            15'd26217: log10_cal = 16'b0000010110100010;
            15'd26218: log10_cal = 16'b0000010110100010;
            15'd26219: log10_cal = 16'b0000010110100010;
            15'd26220: log10_cal = 16'b0000010110100010;
            15'd26221: log10_cal = 16'b0000010110100010;
            15'd26222: log10_cal = 16'b0000010110100010;
            15'd26223: log10_cal = 16'b0000010110100010;
            15'd26224: log10_cal = 16'b0000010110100010;
            15'd26225: log10_cal = 16'b0000010110100010;
            15'd26226: log10_cal = 16'b0000010110100010;
            15'd26227: log10_cal = 16'b0000010110100010;
            15'd26228: log10_cal = 16'b0000010110100010;
            15'd26229: log10_cal = 16'b0000010110100010;
            15'd26230: log10_cal = 16'b0000010110100010;
            15'd26231: log10_cal = 16'b0000010110100010;
            15'd26232: log10_cal = 16'b0000010110100010;
            15'd26233: log10_cal = 16'b0000010110100010;
            15'd26234: log10_cal = 16'b0000010110100010;
            15'd26235: log10_cal = 16'b0000010110100010;
            15'd26236: log10_cal = 16'b0000010110100010;
            15'd26237: log10_cal = 16'b0000010110100010;
            15'd26238: log10_cal = 16'b0000010110100010;
            15'd26239: log10_cal = 16'b0000010110100010;
            15'd26240: log10_cal = 16'b0000010110100010;
            15'd26241: log10_cal = 16'b0000010110100010;
            15'd26242: log10_cal = 16'b0000010110100010;
            15'd26243: log10_cal = 16'b0000010110100010;
            15'd26244: log10_cal = 16'b0000010110100010;
            15'd26245: log10_cal = 16'b0000010110100010;
            15'd26246: log10_cal = 16'b0000010110100010;
            15'd26247: log10_cal = 16'b0000010110100010;
            15'd26248: log10_cal = 16'b0000010110100010;
            15'd26249: log10_cal = 16'b0000010110100010;
            15'd26250: log10_cal = 16'b0000010110100010;
            15'd26251: log10_cal = 16'b0000010110100010;
            15'd26252: log10_cal = 16'b0000010110100010;
            15'd26253: log10_cal = 16'b0000010110100010;
            15'd26254: log10_cal = 16'b0000010110100010;
            15'd26255: log10_cal = 16'b0000010110100010;
            15'd26256: log10_cal = 16'b0000010110100010;
            15'd26257: log10_cal = 16'b0000010110100010;
            15'd26258: log10_cal = 16'b0000010110100010;
            15'd26259: log10_cal = 16'b0000010110100010;
            15'd26260: log10_cal = 16'b0000010110100010;
            15'd26261: log10_cal = 16'b0000010110100010;
            15'd26262: log10_cal = 16'b0000010110100010;
            15'd26263: log10_cal = 16'b0000010110100010;
            15'd26264: log10_cal = 16'b0000010110100010;
            15'd26265: log10_cal = 16'b0000010110100010;
            15'd26266: log10_cal = 16'b0000010110100010;
            15'd26267: log10_cal = 16'b0000010110100010;
            15'd26268: log10_cal = 16'b0000010110100010;
            15'd26269: log10_cal = 16'b0000010110100010;
            15'd26270: log10_cal = 16'b0000010110100010;
            15'd26271: log10_cal = 16'b0000010110100010;
            15'd26272: log10_cal = 16'b0000010110100011;
            15'd26273: log10_cal = 16'b0000010110100011;
            15'd26274: log10_cal = 16'b0000010110100011;
            15'd26275: log10_cal = 16'b0000010110100011;
            15'd26276: log10_cal = 16'b0000010110100011;
            15'd26277: log10_cal = 16'b0000010110100011;
            15'd26278: log10_cal = 16'b0000010110100011;
            15'd26279: log10_cal = 16'b0000010110100011;
            15'd26280: log10_cal = 16'b0000010110100011;
            15'd26281: log10_cal = 16'b0000010110100011;
            15'd26282: log10_cal = 16'b0000010110100011;
            15'd26283: log10_cal = 16'b0000010110100011;
            15'd26284: log10_cal = 16'b0000010110100011;
            15'd26285: log10_cal = 16'b0000010110100011;
            15'd26286: log10_cal = 16'b0000010110100011;
            15'd26287: log10_cal = 16'b0000010110100011;
            15'd26288: log10_cal = 16'b0000010110100011;
            15'd26289: log10_cal = 16'b0000010110100011;
            15'd26290: log10_cal = 16'b0000010110100011;
            15'd26291: log10_cal = 16'b0000010110100011;
            15'd26292: log10_cal = 16'b0000010110100011;
            15'd26293: log10_cal = 16'b0000010110100011;
            15'd26294: log10_cal = 16'b0000010110100011;
            15'd26295: log10_cal = 16'b0000010110100011;
            15'd26296: log10_cal = 16'b0000010110100011;
            15'd26297: log10_cal = 16'b0000010110100011;
            15'd26298: log10_cal = 16'b0000010110100011;
            15'd26299: log10_cal = 16'b0000010110100011;
            15'd26300: log10_cal = 16'b0000010110100011;
            15'd26301: log10_cal = 16'b0000010110100011;
            15'd26302: log10_cal = 16'b0000010110100011;
            15'd26303: log10_cal = 16'b0000010110100011;
            15'd26304: log10_cal = 16'b0000010110100011;
            15'd26305: log10_cal = 16'b0000010110100011;
            15'd26306: log10_cal = 16'b0000010110100011;
            15'd26307: log10_cal = 16'b0000010110100011;
            15'd26308: log10_cal = 16'b0000010110100011;
            15'd26309: log10_cal = 16'b0000010110100011;
            15'd26310: log10_cal = 16'b0000010110100011;
            15'd26311: log10_cal = 16'b0000010110100011;
            15'd26312: log10_cal = 16'b0000010110100011;
            15'd26313: log10_cal = 16'b0000010110100011;
            15'd26314: log10_cal = 16'b0000010110100011;
            15'd26315: log10_cal = 16'b0000010110100011;
            15'd26316: log10_cal = 16'b0000010110100011;
            15'd26317: log10_cal = 16'b0000010110100011;
            15'd26318: log10_cal = 16'b0000010110100011;
            15'd26319: log10_cal = 16'b0000010110100011;
            15'd26320: log10_cal = 16'b0000010110100011;
            15'd26321: log10_cal = 16'b0000010110100011;
            15'd26322: log10_cal = 16'b0000010110100011;
            15'd26323: log10_cal = 16'b0000010110100011;
            15'd26324: log10_cal = 16'b0000010110100011;
            15'd26325: log10_cal = 16'b0000010110100011;
            15'd26326: log10_cal = 16'b0000010110100011;
            15'd26327: log10_cal = 16'b0000010110100011;
            15'd26328: log10_cal = 16'b0000010110100011;
            15'd26329: log10_cal = 16'b0000010110100011;
            15'd26330: log10_cal = 16'b0000010110100011;
            15'd26331: log10_cal = 16'b0000010110100100;
            15'd26332: log10_cal = 16'b0000010110100100;
            15'd26333: log10_cal = 16'b0000010110100100;
            15'd26334: log10_cal = 16'b0000010110100100;
            15'd26335: log10_cal = 16'b0000010110100100;
            15'd26336: log10_cal = 16'b0000010110100100;
            15'd26337: log10_cal = 16'b0000010110100100;
            15'd26338: log10_cal = 16'b0000010110100100;
            15'd26339: log10_cal = 16'b0000010110100100;
            15'd26340: log10_cal = 16'b0000010110100100;
            15'd26341: log10_cal = 16'b0000010110100100;
            15'd26342: log10_cal = 16'b0000010110100100;
            15'd26343: log10_cal = 16'b0000010110100100;
            15'd26344: log10_cal = 16'b0000010110100100;
            15'd26345: log10_cal = 16'b0000010110100100;
            15'd26346: log10_cal = 16'b0000010110100100;
            15'd26347: log10_cal = 16'b0000010110100100;
            15'd26348: log10_cal = 16'b0000010110100100;
            15'd26349: log10_cal = 16'b0000010110100100;
            15'd26350: log10_cal = 16'b0000010110100100;
            15'd26351: log10_cal = 16'b0000010110100100;
            15'd26352: log10_cal = 16'b0000010110100100;
            15'd26353: log10_cal = 16'b0000010110100100;
            15'd26354: log10_cal = 16'b0000010110100100;
            15'd26355: log10_cal = 16'b0000010110100100;
            15'd26356: log10_cal = 16'b0000010110100100;
            15'd26357: log10_cal = 16'b0000010110100100;
            15'd26358: log10_cal = 16'b0000010110100100;
            15'd26359: log10_cal = 16'b0000010110100100;
            15'd26360: log10_cal = 16'b0000010110100100;
            15'd26361: log10_cal = 16'b0000010110100100;
            15'd26362: log10_cal = 16'b0000010110100100;
            15'd26363: log10_cal = 16'b0000010110100100;
            15'd26364: log10_cal = 16'b0000010110100100;
            15'd26365: log10_cal = 16'b0000010110100100;
            15'd26366: log10_cal = 16'b0000010110100100;
            15'd26367: log10_cal = 16'b0000010110100100;
            15'd26368: log10_cal = 16'b0000010110100100;
            15'd26369: log10_cal = 16'b0000010110100100;
            15'd26370: log10_cal = 16'b0000010110100100;
            15'd26371: log10_cal = 16'b0000010110100100;
            15'd26372: log10_cal = 16'b0000010110100100;
            15'd26373: log10_cal = 16'b0000010110100100;
            15'd26374: log10_cal = 16'b0000010110100100;
            15'd26375: log10_cal = 16'b0000010110100100;
            15'd26376: log10_cal = 16'b0000010110100100;
            15'd26377: log10_cal = 16'b0000010110100100;
            15'd26378: log10_cal = 16'b0000010110100100;
            15'd26379: log10_cal = 16'b0000010110100100;
            15'd26380: log10_cal = 16'b0000010110100100;
            15'd26381: log10_cal = 16'b0000010110100100;
            15'd26382: log10_cal = 16'b0000010110100100;
            15'd26383: log10_cal = 16'b0000010110100100;
            15'd26384: log10_cal = 16'b0000010110100100;
            15'd26385: log10_cal = 16'b0000010110100100;
            15'd26386: log10_cal = 16'b0000010110100100;
            15'd26387: log10_cal = 16'b0000010110100100;
            15'd26388: log10_cal = 16'b0000010110100100;
            15'd26389: log10_cal = 16'b0000010110100100;
            15'd26390: log10_cal = 16'b0000010110100101;
            15'd26391: log10_cal = 16'b0000010110100101;
            15'd26392: log10_cal = 16'b0000010110100101;
            15'd26393: log10_cal = 16'b0000010110100101;
            15'd26394: log10_cal = 16'b0000010110100101;
            15'd26395: log10_cal = 16'b0000010110100101;
            15'd26396: log10_cal = 16'b0000010110100101;
            15'd26397: log10_cal = 16'b0000010110100101;
            15'd26398: log10_cal = 16'b0000010110100101;
            15'd26399: log10_cal = 16'b0000010110100101;
            15'd26400: log10_cal = 16'b0000010110100101;
            15'd26401: log10_cal = 16'b0000010110100101;
            15'd26402: log10_cal = 16'b0000010110100101;
            15'd26403: log10_cal = 16'b0000010110100101;
            15'd26404: log10_cal = 16'b0000010110100101;
            15'd26405: log10_cal = 16'b0000010110100101;
            15'd26406: log10_cal = 16'b0000010110100101;
            15'd26407: log10_cal = 16'b0000010110100101;
            15'd26408: log10_cal = 16'b0000010110100101;
            15'd26409: log10_cal = 16'b0000010110100101;
            15'd26410: log10_cal = 16'b0000010110100101;
            15'd26411: log10_cal = 16'b0000010110100101;
            15'd26412: log10_cal = 16'b0000010110100101;
            15'd26413: log10_cal = 16'b0000010110100101;
            15'd26414: log10_cal = 16'b0000010110100101;
            15'd26415: log10_cal = 16'b0000010110100101;
            15'd26416: log10_cal = 16'b0000010110100101;
            15'd26417: log10_cal = 16'b0000010110100101;
            15'd26418: log10_cal = 16'b0000010110100101;
            15'd26419: log10_cal = 16'b0000010110100101;
            15'd26420: log10_cal = 16'b0000010110100101;
            15'd26421: log10_cal = 16'b0000010110100101;
            15'd26422: log10_cal = 16'b0000010110100101;
            15'd26423: log10_cal = 16'b0000010110100101;
            15'd26424: log10_cal = 16'b0000010110100101;
            15'd26425: log10_cal = 16'b0000010110100101;
            15'd26426: log10_cal = 16'b0000010110100101;
            15'd26427: log10_cal = 16'b0000010110100101;
            15'd26428: log10_cal = 16'b0000010110100101;
            15'd26429: log10_cal = 16'b0000010110100101;
            15'd26430: log10_cal = 16'b0000010110100101;
            15'd26431: log10_cal = 16'b0000010110100101;
            15'd26432: log10_cal = 16'b0000010110100101;
            15'd26433: log10_cal = 16'b0000010110100101;
            15'd26434: log10_cal = 16'b0000010110100101;
            15'd26435: log10_cal = 16'b0000010110100101;
            15'd26436: log10_cal = 16'b0000010110100101;
            15'd26437: log10_cal = 16'b0000010110100101;
            15'd26438: log10_cal = 16'b0000010110100101;
            15'd26439: log10_cal = 16'b0000010110100101;
            15'd26440: log10_cal = 16'b0000010110100101;
            15'd26441: log10_cal = 16'b0000010110100101;
            15'd26442: log10_cal = 16'b0000010110100101;
            15'd26443: log10_cal = 16'b0000010110100101;
            15'd26444: log10_cal = 16'b0000010110100101;
            15'd26445: log10_cal = 16'b0000010110100101;
            15'd26446: log10_cal = 16'b0000010110100101;
            15'd26447: log10_cal = 16'b0000010110100101;
            15'd26448: log10_cal = 16'b0000010110100101;
            15'd26449: log10_cal = 16'b0000010110100101;
            15'd26450: log10_cal = 16'b0000010110100110;
            15'd26451: log10_cal = 16'b0000010110100110;
            15'd26452: log10_cal = 16'b0000010110100110;
            15'd26453: log10_cal = 16'b0000010110100110;
            15'd26454: log10_cal = 16'b0000010110100110;
            15'd26455: log10_cal = 16'b0000010110100110;
            15'd26456: log10_cal = 16'b0000010110100110;
            15'd26457: log10_cal = 16'b0000010110100110;
            15'd26458: log10_cal = 16'b0000010110100110;
            15'd26459: log10_cal = 16'b0000010110100110;
            15'd26460: log10_cal = 16'b0000010110100110;
            15'd26461: log10_cal = 16'b0000010110100110;
            15'd26462: log10_cal = 16'b0000010110100110;
            15'd26463: log10_cal = 16'b0000010110100110;
            15'd26464: log10_cal = 16'b0000010110100110;
            15'd26465: log10_cal = 16'b0000010110100110;
            15'd26466: log10_cal = 16'b0000010110100110;
            15'd26467: log10_cal = 16'b0000010110100110;
            15'd26468: log10_cal = 16'b0000010110100110;
            15'd26469: log10_cal = 16'b0000010110100110;
            15'd26470: log10_cal = 16'b0000010110100110;
            15'd26471: log10_cal = 16'b0000010110100110;
            15'd26472: log10_cal = 16'b0000010110100110;
            15'd26473: log10_cal = 16'b0000010110100110;
            15'd26474: log10_cal = 16'b0000010110100110;
            15'd26475: log10_cal = 16'b0000010110100110;
            15'd26476: log10_cal = 16'b0000010110100110;
            15'd26477: log10_cal = 16'b0000010110100110;
            15'd26478: log10_cal = 16'b0000010110100110;
            15'd26479: log10_cal = 16'b0000010110100110;
            15'd26480: log10_cal = 16'b0000010110100110;
            15'd26481: log10_cal = 16'b0000010110100110;
            15'd26482: log10_cal = 16'b0000010110100110;
            15'd26483: log10_cal = 16'b0000010110100110;
            15'd26484: log10_cal = 16'b0000010110100110;
            15'd26485: log10_cal = 16'b0000010110100110;
            15'd26486: log10_cal = 16'b0000010110100110;
            15'd26487: log10_cal = 16'b0000010110100110;
            15'd26488: log10_cal = 16'b0000010110100110;
            15'd26489: log10_cal = 16'b0000010110100110;
            15'd26490: log10_cal = 16'b0000010110100110;
            15'd26491: log10_cal = 16'b0000010110100110;
            15'd26492: log10_cal = 16'b0000010110100110;
            15'd26493: log10_cal = 16'b0000010110100110;
            15'd26494: log10_cal = 16'b0000010110100110;
            15'd26495: log10_cal = 16'b0000010110100110;
            15'd26496: log10_cal = 16'b0000010110100110;
            15'd26497: log10_cal = 16'b0000010110100110;
            15'd26498: log10_cal = 16'b0000010110100110;
            15'd26499: log10_cal = 16'b0000010110100110;
            15'd26500: log10_cal = 16'b0000010110100110;
            15'd26501: log10_cal = 16'b0000010110100110;
            15'd26502: log10_cal = 16'b0000010110100110;
            15'd26503: log10_cal = 16'b0000010110100110;
            15'd26504: log10_cal = 16'b0000010110100110;
            15'd26505: log10_cal = 16'b0000010110100110;
            15'd26506: log10_cal = 16'b0000010110100110;
            15'd26507: log10_cal = 16'b0000010110100110;
            15'd26508: log10_cal = 16'b0000010110100110;
            15'd26509: log10_cal = 16'b0000010110100111;
            15'd26510: log10_cal = 16'b0000010110100111;
            15'd26511: log10_cal = 16'b0000010110100111;
            15'd26512: log10_cal = 16'b0000010110100111;
            15'd26513: log10_cal = 16'b0000010110100111;
            15'd26514: log10_cal = 16'b0000010110100111;
            15'd26515: log10_cal = 16'b0000010110100111;
            15'd26516: log10_cal = 16'b0000010110100111;
            15'd26517: log10_cal = 16'b0000010110100111;
            15'd26518: log10_cal = 16'b0000010110100111;
            15'd26519: log10_cal = 16'b0000010110100111;
            15'd26520: log10_cal = 16'b0000010110100111;
            15'd26521: log10_cal = 16'b0000010110100111;
            15'd26522: log10_cal = 16'b0000010110100111;
            15'd26523: log10_cal = 16'b0000010110100111;
            15'd26524: log10_cal = 16'b0000010110100111;
            15'd26525: log10_cal = 16'b0000010110100111;
            15'd26526: log10_cal = 16'b0000010110100111;
            15'd26527: log10_cal = 16'b0000010110100111;
            15'd26528: log10_cal = 16'b0000010110100111;
            15'd26529: log10_cal = 16'b0000010110100111;
            15'd26530: log10_cal = 16'b0000010110100111;
            15'd26531: log10_cal = 16'b0000010110100111;
            15'd26532: log10_cal = 16'b0000010110100111;
            15'd26533: log10_cal = 16'b0000010110100111;
            15'd26534: log10_cal = 16'b0000010110100111;
            15'd26535: log10_cal = 16'b0000010110100111;
            15'd26536: log10_cal = 16'b0000010110100111;
            15'd26537: log10_cal = 16'b0000010110100111;
            15'd26538: log10_cal = 16'b0000010110100111;
            15'd26539: log10_cal = 16'b0000010110100111;
            15'd26540: log10_cal = 16'b0000010110100111;
            15'd26541: log10_cal = 16'b0000010110100111;
            15'd26542: log10_cal = 16'b0000010110100111;
            15'd26543: log10_cal = 16'b0000010110100111;
            15'd26544: log10_cal = 16'b0000010110100111;
            15'd26545: log10_cal = 16'b0000010110100111;
            15'd26546: log10_cal = 16'b0000010110100111;
            15'd26547: log10_cal = 16'b0000010110100111;
            15'd26548: log10_cal = 16'b0000010110100111;
            15'd26549: log10_cal = 16'b0000010110100111;
            15'd26550: log10_cal = 16'b0000010110100111;
            15'd26551: log10_cal = 16'b0000010110100111;
            15'd26552: log10_cal = 16'b0000010110100111;
            15'd26553: log10_cal = 16'b0000010110100111;
            15'd26554: log10_cal = 16'b0000010110100111;
            15'd26555: log10_cal = 16'b0000010110100111;
            15'd26556: log10_cal = 16'b0000010110100111;
            15'd26557: log10_cal = 16'b0000010110100111;
            15'd26558: log10_cal = 16'b0000010110100111;
            15'd26559: log10_cal = 16'b0000010110100111;
            15'd26560: log10_cal = 16'b0000010110100111;
            15'd26561: log10_cal = 16'b0000010110100111;
            15'd26562: log10_cal = 16'b0000010110100111;
            15'd26563: log10_cal = 16'b0000010110100111;
            15'd26564: log10_cal = 16'b0000010110100111;
            15'd26565: log10_cal = 16'b0000010110100111;
            15'd26566: log10_cal = 16'b0000010110100111;
            15'd26567: log10_cal = 16'b0000010110100111;
            15'd26568: log10_cal = 16'b0000010110100111;
            15'd26569: log10_cal = 16'b0000010110101000;
            15'd26570: log10_cal = 16'b0000010110101000;
            15'd26571: log10_cal = 16'b0000010110101000;
            15'd26572: log10_cal = 16'b0000010110101000;
            15'd26573: log10_cal = 16'b0000010110101000;
            15'd26574: log10_cal = 16'b0000010110101000;
            15'd26575: log10_cal = 16'b0000010110101000;
            15'd26576: log10_cal = 16'b0000010110101000;
            15'd26577: log10_cal = 16'b0000010110101000;
            15'd26578: log10_cal = 16'b0000010110101000;
            15'd26579: log10_cal = 16'b0000010110101000;
            15'd26580: log10_cal = 16'b0000010110101000;
            15'd26581: log10_cal = 16'b0000010110101000;
            15'd26582: log10_cal = 16'b0000010110101000;
            15'd26583: log10_cal = 16'b0000010110101000;
            15'd26584: log10_cal = 16'b0000010110101000;
            15'd26585: log10_cal = 16'b0000010110101000;
            15'd26586: log10_cal = 16'b0000010110101000;
            15'd26587: log10_cal = 16'b0000010110101000;
            15'd26588: log10_cal = 16'b0000010110101000;
            15'd26589: log10_cal = 16'b0000010110101000;
            15'd26590: log10_cal = 16'b0000010110101000;
            15'd26591: log10_cal = 16'b0000010110101000;
            15'd26592: log10_cal = 16'b0000010110101000;
            15'd26593: log10_cal = 16'b0000010110101000;
            15'd26594: log10_cal = 16'b0000010110101000;
            15'd26595: log10_cal = 16'b0000010110101000;
            15'd26596: log10_cal = 16'b0000010110101000;
            15'd26597: log10_cal = 16'b0000010110101000;
            15'd26598: log10_cal = 16'b0000010110101000;
            15'd26599: log10_cal = 16'b0000010110101000;
            15'd26600: log10_cal = 16'b0000010110101000;
            15'd26601: log10_cal = 16'b0000010110101000;
            15'd26602: log10_cal = 16'b0000010110101000;
            15'd26603: log10_cal = 16'b0000010110101000;
            15'd26604: log10_cal = 16'b0000010110101000;
            15'd26605: log10_cal = 16'b0000010110101000;
            15'd26606: log10_cal = 16'b0000010110101000;
            15'd26607: log10_cal = 16'b0000010110101000;
            15'd26608: log10_cal = 16'b0000010110101000;
            15'd26609: log10_cal = 16'b0000010110101000;
            15'd26610: log10_cal = 16'b0000010110101000;
            15'd26611: log10_cal = 16'b0000010110101000;
            15'd26612: log10_cal = 16'b0000010110101000;
            15'd26613: log10_cal = 16'b0000010110101000;
            15'd26614: log10_cal = 16'b0000010110101000;
            15'd26615: log10_cal = 16'b0000010110101000;
            15'd26616: log10_cal = 16'b0000010110101000;
            15'd26617: log10_cal = 16'b0000010110101000;
            15'd26618: log10_cal = 16'b0000010110101000;
            15'd26619: log10_cal = 16'b0000010110101000;
            15'd26620: log10_cal = 16'b0000010110101000;
            15'd26621: log10_cal = 16'b0000010110101000;
            15'd26622: log10_cal = 16'b0000010110101000;
            15'd26623: log10_cal = 16'b0000010110101000;
            15'd26624: log10_cal = 16'b0000010110101000;
            15'd26625: log10_cal = 16'b0000010110101000;
            15'd26626: log10_cal = 16'b0000010110101000;
            15'd26627: log10_cal = 16'b0000010110101000;
            15'd26628: log10_cal = 16'b0000010110101000;
            15'd26629: log10_cal = 16'b0000010110101001;
            15'd26630: log10_cal = 16'b0000010110101001;
            15'd26631: log10_cal = 16'b0000010110101001;
            15'd26632: log10_cal = 16'b0000010110101001;
            15'd26633: log10_cal = 16'b0000010110101001;
            15'd26634: log10_cal = 16'b0000010110101001;
            15'd26635: log10_cal = 16'b0000010110101001;
            15'd26636: log10_cal = 16'b0000010110101001;
            15'd26637: log10_cal = 16'b0000010110101001;
            15'd26638: log10_cal = 16'b0000010110101001;
            15'd26639: log10_cal = 16'b0000010110101001;
            15'd26640: log10_cal = 16'b0000010110101001;
            15'd26641: log10_cal = 16'b0000010110101001;
            15'd26642: log10_cal = 16'b0000010110101001;
            15'd26643: log10_cal = 16'b0000010110101001;
            15'd26644: log10_cal = 16'b0000010110101001;
            15'd26645: log10_cal = 16'b0000010110101001;
            15'd26646: log10_cal = 16'b0000010110101001;
            15'd26647: log10_cal = 16'b0000010110101001;
            15'd26648: log10_cal = 16'b0000010110101001;
            15'd26649: log10_cal = 16'b0000010110101001;
            15'd26650: log10_cal = 16'b0000010110101001;
            15'd26651: log10_cal = 16'b0000010110101001;
            15'd26652: log10_cal = 16'b0000010110101001;
            15'd26653: log10_cal = 16'b0000010110101001;
            15'd26654: log10_cal = 16'b0000010110101001;
            15'd26655: log10_cal = 16'b0000010110101001;
            15'd26656: log10_cal = 16'b0000010110101001;
            15'd26657: log10_cal = 16'b0000010110101001;
            15'd26658: log10_cal = 16'b0000010110101001;
            15'd26659: log10_cal = 16'b0000010110101001;
            15'd26660: log10_cal = 16'b0000010110101001;
            15'd26661: log10_cal = 16'b0000010110101001;
            15'd26662: log10_cal = 16'b0000010110101001;
            15'd26663: log10_cal = 16'b0000010110101001;
            15'd26664: log10_cal = 16'b0000010110101001;
            15'd26665: log10_cal = 16'b0000010110101001;
            15'd26666: log10_cal = 16'b0000010110101001;
            15'd26667: log10_cal = 16'b0000010110101001;
            15'd26668: log10_cal = 16'b0000010110101001;
            15'd26669: log10_cal = 16'b0000010110101001;
            15'd26670: log10_cal = 16'b0000010110101001;
            15'd26671: log10_cal = 16'b0000010110101001;
            15'd26672: log10_cal = 16'b0000010110101001;
            15'd26673: log10_cal = 16'b0000010110101001;
            15'd26674: log10_cal = 16'b0000010110101001;
            15'd26675: log10_cal = 16'b0000010110101001;
            15'd26676: log10_cal = 16'b0000010110101001;
            15'd26677: log10_cal = 16'b0000010110101001;
            15'd26678: log10_cal = 16'b0000010110101001;
            15'd26679: log10_cal = 16'b0000010110101001;
            15'd26680: log10_cal = 16'b0000010110101001;
            15'd26681: log10_cal = 16'b0000010110101001;
            15'd26682: log10_cal = 16'b0000010110101001;
            15'd26683: log10_cal = 16'b0000010110101001;
            15'd26684: log10_cal = 16'b0000010110101001;
            15'd26685: log10_cal = 16'b0000010110101001;
            15'd26686: log10_cal = 16'b0000010110101001;
            15'd26687: log10_cal = 16'b0000010110101001;
            15'd26688: log10_cal = 16'b0000010110101010;
            15'd26689: log10_cal = 16'b0000010110101010;
            15'd26690: log10_cal = 16'b0000010110101010;
            15'd26691: log10_cal = 16'b0000010110101010;
            15'd26692: log10_cal = 16'b0000010110101010;
            15'd26693: log10_cal = 16'b0000010110101010;
            15'd26694: log10_cal = 16'b0000010110101010;
            15'd26695: log10_cal = 16'b0000010110101010;
            15'd26696: log10_cal = 16'b0000010110101010;
            15'd26697: log10_cal = 16'b0000010110101010;
            15'd26698: log10_cal = 16'b0000010110101010;
            15'd26699: log10_cal = 16'b0000010110101010;
            15'd26700: log10_cal = 16'b0000010110101010;
            15'd26701: log10_cal = 16'b0000010110101010;
            15'd26702: log10_cal = 16'b0000010110101010;
            15'd26703: log10_cal = 16'b0000010110101010;
            15'd26704: log10_cal = 16'b0000010110101010;
            15'd26705: log10_cal = 16'b0000010110101010;
            15'd26706: log10_cal = 16'b0000010110101010;
            15'd26707: log10_cal = 16'b0000010110101010;
            15'd26708: log10_cal = 16'b0000010110101010;
            15'd26709: log10_cal = 16'b0000010110101010;
            15'd26710: log10_cal = 16'b0000010110101010;
            15'd26711: log10_cal = 16'b0000010110101010;
            15'd26712: log10_cal = 16'b0000010110101010;
            15'd26713: log10_cal = 16'b0000010110101010;
            15'd26714: log10_cal = 16'b0000010110101010;
            15'd26715: log10_cal = 16'b0000010110101010;
            15'd26716: log10_cal = 16'b0000010110101010;
            15'd26717: log10_cal = 16'b0000010110101010;
            15'd26718: log10_cal = 16'b0000010110101010;
            15'd26719: log10_cal = 16'b0000010110101010;
            15'd26720: log10_cal = 16'b0000010110101010;
            15'd26721: log10_cal = 16'b0000010110101010;
            15'd26722: log10_cal = 16'b0000010110101010;
            15'd26723: log10_cal = 16'b0000010110101010;
            15'd26724: log10_cal = 16'b0000010110101010;
            15'd26725: log10_cal = 16'b0000010110101010;
            15'd26726: log10_cal = 16'b0000010110101010;
            15'd26727: log10_cal = 16'b0000010110101010;
            15'd26728: log10_cal = 16'b0000010110101010;
            15'd26729: log10_cal = 16'b0000010110101010;
            15'd26730: log10_cal = 16'b0000010110101010;
            15'd26731: log10_cal = 16'b0000010110101010;
            15'd26732: log10_cal = 16'b0000010110101010;
            15'd26733: log10_cal = 16'b0000010110101010;
            15'd26734: log10_cal = 16'b0000010110101010;
            15'd26735: log10_cal = 16'b0000010110101010;
            15'd26736: log10_cal = 16'b0000010110101010;
            15'd26737: log10_cal = 16'b0000010110101010;
            15'd26738: log10_cal = 16'b0000010110101010;
            15'd26739: log10_cal = 16'b0000010110101010;
            15'd26740: log10_cal = 16'b0000010110101010;
            15'd26741: log10_cal = 16'b0000010110101010;
            15'd26742: log10_cal = 16'b0000010110101010;
            15'd26743: log10_cal = 16'b0000010110101010;
            15'd26744: log10_cal = 16'b0000010110101010;
            15'd26745: log10_cal = 16'b0000010110101010;
            15'd26746: log10_cal = 16'b0000010110101010;
            15'd26747: log10_cal = 16'b0000010110101010;
            15'd26748: log10_cal = 16'b0000010110101010;
            15'd26749: log10_cal = 16'b0000010110101011;
            15'd26750: log10_cal = 16'b0000010110101011;
            15'd26751: log10_cal = 16'b0000010110101011;
            15'd26752: log10_cal = 16'b0000010110101011;
            15'd26753: log10_cal = 16'b0000010110101011;
            15'd26754: log10_cal = 16'b0000010110101011;
            15'd26755: log10_cal = 16'b0000010110101011;
            15'd26756: log10_cal = 16'b0000010110101011;
            15'd26757: log10_cal = 16'b0000010110101011;
            15'd26758: log10_cal = 16'b0000010110101011;
            15'd26759: log10_cal = 16'b0000010110101011;
            15'd26760: log10_cal = 16'b0000010110101011;
            15'd26761: log10_cal = 16'b0000010110101011;
            15'd26762: log10_cal = 16'b0000010110101011;
            15'd26763: log10_cal = 16'b0000010110101011;
            15'd26764: log10_cal = 16'b0000010110101011;
            15'd26765: log10_cal = 16'b0000010110101011;
            15'd26766: log10_cal = 16'b0000010110101011;
            15'd26767: log10_cal = 16'b0000010110101011;
            15'd26768: log10_cal = 16'b0000010110101011;
            15'd26769: log10_cal = 16'b0000010110101011;
            15'd26770: log10_cal = 16'b0000010110101011;
            15'd26771: log10_cal = 16'b0000010110101011;
            15'd26772: log10_cal = 16'b0000010110101011;
            15'd26773: log10_cal = 16'b0000010110101011;
            15'd26774: log10_cal = 16'b0000010110101011;
            15'd26775: log10_cal = 16'b0000010110101011;
            15'd26776: log10_cal = 16'b0000010110101011;
            15'd26777: log10_cal = 16'b0000010110101011;
            15'd26778: log10_cal = 16'b0000010110101011;
            15'd26779: log10_cal = 16'b0000010110101011;
            15'd26780: log10_cal = 16'b0000010110101011;
            15'd26781: log10_cal = 16'b0000010110101011;
            15'd26782: log10_cal = 16'b0000010110101011;
            15'd26783: log10_cal = 16'b0000010110101011;
            15'd26784: log10_cal = 16'b0000010110101011;
            15'd26785: log10_cal = 16'b0000010110101011;
            15'd26786: log10_cal = 16'b0000010110101011;
            15'd26787: log10_cal = 16'b0000010110101011;
            15'd26788: log10_cal = 16'b0000010110101011;
            15'd26789: log10_cal = 16'b0000010110101011;
            15'd26790: log10_cal = 16'b0000010110101011;
            15'd26791: log10_cal = 16'b0000010110101011;
            15'd26792: log10_cal = 16'b0000010110101011;
            15'd26793: log10_cal = 16'b0000010110101011;
            15'd26794: log10_cal = 16'b0000010110101011;
            15'd26795: log10_cal = 16'b0000010110101011;
            15'd26796: log10_cal = 16'b0000010110101011;
            15'd26797: log10_cal = 16'b0000010110101011;
            15'd26798: log10_cal = 16'b0000010110101011;
            15'd26799: log10_cal = 16'b0000010110101011;
            15'd26800: log10_cal = 16'b0000010110101011;
            15'd26801: log10_cal = 16'b0000010110101011;
            15'd26802: log10_cal = 16'b0000010110101011;
            15'd26803: log10_cal = 16'b0000010110101011;
            15'd26804: log10_cal = 16'b0000010110101011;
            15'd26805: log10_cal = 16'b0000010110101011;
            15'd26806: log10_cal = 16'b0000010110101011;
            15'd26807: log10_cal = 16'b0000010110101011;
            15'd26808: log10_cal = 16'b0000010110101011;
            15'd26809: log10_cal = 16'b0000010110101100;
            15'd26810: log10_cal = 16'b0000010110101100;
            15'd26811: log10_cal = 16'b0000010110101100;
            15'd26812: log10_cal = 16'b0000010110101100;
            15'd26813: log10_cal = 16'b0000010110101100;
            15'd26814: log10_cal = 16'b0000010110101100;
            15'd26815: log10_cal = 16'b0000010110101100;
            15'd26816: log10_cal = 16'b0000010110101100;
            15'd26817: log10_cal = 16'b0000010110101100;
            15'd26818: log10_cal = 16'b0000010110101100;
            15'd26819: log10_cal = 16'b0000010110101100;
            15'd26820: log10_cal = 16'b0000010110101100;
            15'd26821: log10_cal = 16'b0000010110101100;
            15'd26822: log10_cal = 16'b0000010110101100;
            15'd26823: log10_cal = 16'b0000010110101100;
            15'd26824: log10_cal = 16'b0000010110101100;
            15'd26825: log10_cal = 16'b0000010110101100;
            15'd26826: log10_cal = 16'b0000010110101100;
            15'd26827: log10_cal = 16'b0000010110101100;
            15'd26828: log10_cal = 16'b0000010110101100;
            15'd26829: log10_cal = 16'b0000010110101100;
            15'd26830: log10_cal = 16'b0000010110101100;
            15'd26831: log10_cal = 16'b0000010110101100;
            15'd26832: log10_cal = 16'b0000010110101100;
            15'd26833: log10_cal = 16'b0000010110101100;
            15'd26834: log10_cal = 16'b0000010110101100;
            15'd26835: log10_cal = 16'b0000010110101100;
            15'd26836: log10_cal = 16'b0000010110101100;
            15'd26837: log10_cal = 16'b0000010110101100;
            15'd26838: log10_cal = 16'b0000010110101100;
            15'd26839: log10_cal = 16'b0000010110101100;
            15'd26840: log10_cal = 16'b0000010110101100;
            15'd26841: log10_cal = 16'b0000010110101100;
            15'd26842: log10_cal = 16'b0000010110101100;
            15'd26843: log10_cal = 16'b0000010110101100;
            15'd26844: log10_cal = 16'b0000010110101100;
            15'd26845: log10_cal = 16'b0000010110101100;
            15'd26846: log10_cal = 16'b0000010110101100;
            15'd26847: log10_cal = 16'b0000010110101100;
            15'd26848: log10_cal = 16'b0000010110101100;
            15'd26849: log10_cal = 16'b0000010110101100;
            15'd26850: log10_cal = 16'b0000010110101100;
            15'd26851: log10_cal = 16'b0000010110101100;
            15'd26852: log10_cal = 16'b0000010110101100;
            15'd26853: log10_cal = 16'b0000010110101100;
            15'd26854: log10_cal = 16'b0000010110101100;
            15'd26855: log10_cal = 16'b0000010110101100;
            15'd26856: log10_cal = 16'b0000010110101100;
            15'd26857: log10_cal = 16'b0000010110101100;
            15'd26858: log10_cal = 16'b0000010110101100;
            15'd26859: log10_cal = 16'b0000010110101100;
            15'd26860: log10_cal = 16'b0000010110101100;
            15'd26861: log10_cal = 16'b0000010110101100;
            15'd26862: log10_cal = 16'b0000010110101100;
            15'd26863: log10_cal = 16'b0000010110101100;
            15'd26864: log10_cal = 16'b0000010110101100;
            15'd26865: log10_cal = 16'b0000010110101100;
            15'd26866: log10_cal = 16'b0000010110101100;
            15'd26867: log10_cal = 16'b0000010110101100;
            15'd26868: log10_cal = 16'b0000010110101100;
            15'd26869: log10_cal = 16'b0000010110101101;
            15'd26870: log10_cal = 16'b0000010110101101;
            15'd26871: log10_cal = 16'b0000010110101101;
            15'd26872: log10_cal = 16'b0000010110101101;
            15'd26873: log10_cal = 16'b0000010110101101;
            15'd26874: log10_cal = 16'b0000010110101101;
            15'd26875: log10_cal = 16'b0000010110101101;
            15'd26876: log10_cal = 16'b0000010110101101;
            15'd26877: log10_cal = 16'b0000010110101101;
            15'd26878: log10_cal = 16'b0000010110101101;
            15'd26879: log10_cal = 16'b0000010110101101;
            15'd26880: log10_cal = 16'b0000010110101101;
            15'd26881: log10_cal = 16'b0000010110101101;
            15'd26882: log10_cal = 16'b0000010110101101;
            15'd26883: log10_cal = 16'b0000010110101101;
            15'd26884: log10_cal = 16'b0000010110101101;
            15'd26885: log10_cal = 16'b0000010110101101;
            15'd26886: log10_cal = 16'b0000010110101101;
            15'd26887: log10_cal = 16'b0000010110101101;
            15'd26888: log10_cal = 16'b0000010110101101;
            15'd26889: log10_cal = 16'b0000010110101101;
            15'd26890: log10_cal = 16'b0000010110101101;
            15'd26891: log10_cal = 16'b0000010110101101;
            15'd26892: log10_cal = 16'b0000010110101101;
            15'd26893: log10_cal = 16'b0000010110101101;
            15'd26894: log10_cal = 16'b0000010110101101;
            15'd26895: log10_cal = 16'b0000010110101101;
            15'd26896: log10_cal = 16'b0000010110101101;
            15'd26897: log10_cal = 16'b0000010110101101;
            15'd26898: log10_cal = 16'b0000010110101101;
            15'd26899: log10_cal = 16'b0000010110101101;
            15'd26900: log10_cal = 16'b0000010110101101;
            15'd26901: log10_cal = 16'b0000010110101101;
            15'd26902: log10_cal = 16'b0000010110101101;
            15'd26903: log10_cal = 16'b0000010110101101;
            15'd26904: log10_cal = 16'b0000010110101101;
            15'd26905: log10_cal = 16'b0000010110101101;
            15'd26906: log10_cal = 16'b0000010110101101;
            15'd26907: log10_cal = 16'b0000010110101101;
            15'd26908: log10_cal = 16'b0000010110101101;
            15'd26909: log10_cal = 16'b0000010110101101;
            15'd26910: log10_cal = 16'b0000010110101101;
            15'd26911: log10_cal = 16'b0000010110101101;
            15'd26912: log10_cal = 16'b0000010110101101;
            15'd26913: log10_cal = 16'b0000010110101101;
            15'd26914: log10_cal = 16'b0000010110101101;
            15'd26915: log10_cal = 16'b0000010110101101;
            15'd26916: log10_cal = 16'b0000010110101101;
            15'd26917: log10_cal = 16'b0000010110101101;
            15'd26918: log10_cal = 16'b0000010110101101;
            15'd26919: log10_cal = 16'b0000010110101101;
            15'd26920: log10_cal = 16'b0000010110101101;
            15'd26921: log10_cal = 16'b0000010110101101;
            15'd26922: log10_cal = 16'b0000010110101101;
            15'd26923: log10_cal = 16'b0000010110101101;
            15'd26924: log10_cal = 16'b0000010110101101;
            15'd26925: log10_cal = 16'b0000010110101101;
            15'd26926: log10_cal = 16'b0000010110101101;
            15'd26927: log10_cal = 16'b0000010110101101;
            15'd26928: log10_cal = 16'b0000010110101101;
            15'd26929: log10_cal = 16'b0000010110101101;
            15'd26930: log10_cal = 16'b0000010110101110;
            15'd26931: log10_cal = 16'b0000010110101110;
            15'd26932: log10_cal = 16'b0000010110101110;
            15'd26933: log10_cal = 16'b0000010110101110;
            15'd26934: log10_cal = 16'b0000010110101110;
            15'd26935: log10_cal = 16'b0000010110101110;
            15'd26936: log10_cal = 16'b0000010110101110;
            15'd26937: log10_cal = 16'b0000010110101110;
            15'd26938: log10_cal = 16'b0000010110101110;
            15'd26939: log10_cal = 16'b0000010110101110;
            15'd26940: log10_cal = 16'b0000010110101110;
            15'd26941: log10_cal = 16'b0000010110101110;
            15'd26942: log10_cal = 16'b0000010110101110;
            15'd26943: log10_cal = 16'b0000010110101110;
            15'd26944: log10_cal = 16'b0000010110101110;
            15'd26945: log10_cal = 16'b0000010110101110;
            15'd26946: log10_cal = 16'b0000010110101110;
            15'd26947: log10_cal = 16'b0000010110101110;
            15'd26948: log10_cal = 16'b0000010110101110;
            15'd26949: log10_cal = 16'b0000010110101110;
            15'd26950: log10_cal = 16'b0000010110101110;
            15'd26951: log10_cal = 16'b0000010110101110;
            15'd26952: log10_cal = 16'b0000010110101110;
            15'd26953: log10_cal = 16'b0000010110101110;
            15'd26954: log10_cal = 16'b0000010110101110;
            15'd26955: log10_cal = 16'b0000010110101110;
            15'd26956: log10_cal = 16'b0000010110101110;
            15'd26957: log10_cal = 16'b0000010110101110;
            15'd26958: log10_cal = 16'b0000010110101110;
            15'd26959: log10_cal = 16'b0000010110101110;
            15'd26960: log10_cal = 16'b0000010110101110;
            15'd26961: log10_cal = 16'b0000010110101110;
            15'd26962: log10_cal = 16'b0000010110101110;
            15'd26963: log10_cal = 16'b0000010110101110;
            15'd26964: log10_cal = 16'b0000010110101110;
            15'd26965: log10_cal = 16'b0000010110101110;
            15'd26966: log10_cal = 16'b0000010110101110;
            15'd26967: log10_cal = 16'b0000010110101110;
            15'd26968: log10_cal = 16'b0000010110101110;
            15'd26969: log10_cal = 16'b0000010110101110;
            15'd26970: log10_cal = 16'b0000010110101110;
            15'd26971: log10_cal = 16'b0000010110101110;
            15'd26972: log10_cal = 16'b0000010110101110;
            15'd26973: log10_cal = 16'b0000010110101110;
            15'd26974: log10_cal = 16'b0000010110101110;
            15'd26975: log10_cal = 16'b0000010110101110;
            15'd26976: log10_cal = 16'b0000010110101110;
            15'd26977: log10_cal = 16'b0000010110101110;
            15'd26978: log10_cal = 16'b0000010110101110;
            15'd26979: log10_cal = 16'b0000010110101110;
            15'd26980: log10_cal = 16'b0000010110101110;
            15'd26981: log10_cal = 16'b0000010110101110;
            15'd26982: log10_cal = 16'b0000010110101110;
            15'd26983: log10_cal = 16'b0000010110101110;
            15'd26984: log10_cal = 16'b0000010110101110;
            15'd26985: log10_cal = 16'b0000010110101110;
            15'd26986: log10_cal = 16'b0000010110101110;
            15'd26987: log10_cal = 16'b0000010110101110;
            15'd26988: log10_cal = 16'b0000010110101110;
            15'd26989: log10_cal = 16'b0000010110101110;
            15'd26990: log10_cal = 16'b0000010110101111;
            15'd26991: log10_cal = 16'b0000010110101111;
            15'd26992: log10_cal = 16'b0000010110101111;
            15'd26993: log10_cal = 16'b0000010110101111;
            15'd26994: log10_cal = 16'b0000010110101111;
            15'd26995: log10_cal = 16'b0000010110101111;
            15'd26996: log10_cal = 16'b0000010110101111;
            15'd26997: log10_cal = 16'b0000010110101111;
            15'd26998: log10_cal = 16'b0000010110101111;
            15'd26999: log10_cal = 16'b0000010110101111;
            15'd27000: log10_cal = 16'b0000010110101111;
            15'd27001: log10_cal = 16'b0000010110101111;
            15'd27002: log10_cal = 16'b0000010110101111;
            15'd27003: log10_cal = 16'b0000010110101111;
            15'd27004: log10_cal = 16'b0000010110101111;
            15'd27005: log10_cal = 16'b0000010110101111;
            15'd27006: log10_cal = 16'b0000010110101111;
            15'd27007: log10_cal = 16'b0000010110101111;
            15'd27008: log10_cal = 16'b0000010110101111;
            15'd27009: log10_cal = 16'b0000010110101111;
            15'd27010: log10_cal = 16'b0000010110101111;
            15'd27011: log10_cal = 16'b0000010110101111;
            15'd27012: log10_cal = 16'b0000010110101111;
            15'd27013: log10_cal = 16'b0000010110101111;
            15'd27014: log10_cal = 16'b0000010110101111;
            15'd27015: log10_cal = 16'b0000010110101111;
            15'd27016: log10_cal = 16'b0000010110101111;
            15'd27017: log10_cal = 16'b0000010110101111;
            15'd27018: log10_cal = 16'b0000010110101111;
            15'd27019: log10_cal = 16'b0000010110101111;
            15'd27020: log10_cal = 16'b0000010110101111;
            15'd27021: log10_cal = 16'b0000010110101111;
            15'd27022: log10_cal = 16'b0000010110101111;
            15'd27023: log10_cal = 16'b0000010110101111;
            15'd27024: log10_cal = 16'b0000010110101111;
            15'd27025: log10_cal = 16'b0000010110101111;
            15'd27026: log10_cal = 16'b0000010110101111;
            15'd27027: log10_cal = 16'b0000010110101111;
            15'd27028: log10_cal = 16'b0000010110101111;
            15'd27029: log10_cal = 16'b0000010110101111;
            15'd27030: log10_cal = 16'b0000010110101111;
            15'd27031: log10_cal = 16'b0000010110101111;
            15'd27032: log10_cal = 16'b0000010110101111;
            15'd27033: log10_cal = 16'b0000010110101111;
            15'd27034: log10_cal = 16'b0000010110101111;
            15'd27035: log10_cal = 16'b0000010110101111;
            15'd27036: log10_cal = 16'b0000010110101111;
            15'd27037: log10_cal = 16'b0000010110101111;
            15'd27038: log10_cal = 16'b0000010110101111;
            15'd27039: log10_cal = 16'b0000010110101111;
            15'd27040: log10_cal = 16'b0000010110101111;
            15'd27041: log10_cal = 16'b0000010110101111;
            15'd27042: log10_cal = 16'b0000010110101111;
            15'd27043: log10_cal = 16'b0000010110101111;
            15'd27044: log10_cal = 16'b0000010110101111;
            15'd27045: log10_cal = 16'b0000010110101111;
            15'd27046: log10_cal = 16'b0000010110101111;
            15'd27047: log10_cal = 16'b0000010110101111;
            15'd27048: log10_cal = 16'b0000010110101111;
            15'd27049: log10_cal = 16'b0000010110101111;
            15'd27050: log10_cal = 16'b0000010110101111;
            15'd27051: log10_cal = 16'b0000010110110000;
            15'd27052: log10_cal = 16'b0000010110110000;
            15'd27053: log10_cal = 16'b0000010110110000;
            15'd27054: log10_cal = 16'b0000010110110000;
            15'd27055: log10_cal = 16'b0000010110110000;
            15'd27056: log10_cal = 16'b0000010110110000;
            15'd27057: log10_cal = 16'b0000010110110000;
            15'd27058: log10_cal = 16'b0000010110110000;
            15'd27059: log10_cal = 16'b0000010110110000;
            15'd27060: log10_cal = 16'b0000010110110000;
            15'd27061: log10_cal = 16'b0000010110110000;
            15'd27062: log10_cal = 16'b0000010110110000;
            15'd27063: log10_cal = 16'b0000010110110000;
            15'd27064: log10_cal = 16'b0000010110110000;
            15'd27065: log10_cal = 16'b0000010110110000;
            15'd27066: log10_cal = 16'b0000010110110000;
            15'd27067: log10_cal = 16'b0000010110110000;
            15'd27068: log10_cal = 16'b0000010110110000;
            15'd27069: log10_cal = 16'b0000010110110000;
            15'd27070: log10_cal = 16'b0000010110110000;
            15'd27071: log10_cal = 16'b0000010110110000;
            15'd27072: log10_cal = 16'b0000010110110000;
            15'd27073: log10_cal = 16'b0000010110110000;
            15'd27074: log10_cal = 16'b0000010110110000;
            15'd27075: log10_cal = 16'b0000010110110000;
            15'd27076: log10_cal = 16'b0000010110110000;
            15'd27077: log10_cal = 16'b0000010110110000;
            15'd27078: log10_cal = 16'b0000010110110000;
            15'd27079: log10_cal = 16'b0000010110110000;
            15'd27080: log10_cal = 16'b0000010110110000;
            15'd27081: log10_cal = 16'b0000010110110000;
            15'd27082: log10_cal = 16'b0000010110110000;
            15'd27083: log10_cal = 16'b0000010110110000;
            15'd27084: log10_cal = 16'b0000010110110000;
            15'd27085: log10_cal = 16'b0000010110110000;
            15'd27086: log10_cal = 16'b0000010110110000;
            15'd27087: log10_cal = 16'b0000010110110000;
            15'd27088: log10_cal = 16'b0000010110110000;
            15'd27089: log10_cal = 16'b0000010110110000;
            15'd27090: log10_cal = 16'b0000010110110000;
            15'd27091: log10_cal = 16'b0000010110110000;
            15'd27092: log10_cal = 16'b0000010110110000;
            15'd27093: log10_cal = 16'b0000010110110000;
            15'd27094: log10_cal = 16'b0000010110110000;
            15'd27095: log10_cal = 16'b0000010110110000;
            15'd27096: log10_cal = 16'b0000010110110000;
            15'd27097: log10_cal = 16'b0000010110110000;
            15'd27098: log10_cal = 16'b0000010110110000;
            15'd27099: log10_cal = 16'b0000010110110000;
            15'd27100: log10_cal = 16'b0000010110110000;
            15'd27101: log10_cal = 16'b0000010110110000;
            15'd27102: log10_cal = 16'b0000010110110000;
            15'd27103: log10_cal = 16'b0000010110110000;
            15'd27104: log10_cal = 16'b0000010110110000;
            15'd27105: log10_cal = 16'b0000010110110000;
            15'd27106: log10_cal = 16'b0000010110110000;
            15'd27107: log10_cal = 16'b0000010110110000;
            15'd27108: log10_cal = 16'b0000010110110000;
            15'd27109: log10_cal = 16'b0000010110110000;
            15'd27110: log10_cal = 16'b0000010110110000;
            15'd27111: log10_cal = 16'b0000010110110000;
            15'd27112: log10_cal = 16'b0000010110110001;
            15'd27113: log10_cal = 16'b0000010110110001;
            15'd27114: log10_cal = 16'b0000010110110001;
            15'd27115: log10_cal = 16'b0000010110110001;
            15'd27116: log10_cal = 16'b0000010110110001;
            15'd27117: log10_cal = 16'b0000010110110001;
            15'd27118: log10_cal = 16'b0000010110110001;
            15'd27119: log10_cal = 16'b0000010110110001;
            15'd27120: log10_cal = 16'b0000010110110001;
            15'd27121: log10_cal = 16'b0000010110110001;
            15'd27122: log10_cal = 16'b0000010110110001;
            15'd27123: log10_cal = 16'b0000010110110001;
            15'd27124: log10_cal = 16'b0000010110110001;
            15'd27125: log10_cal = 16'b0000010110110001;
            15'd27126: log10_cal = 16'b0000010110110001;
            15'd27127: log10_cal = 16'b0000010110110001;
            15'd27128: log10_cal = 16'b0000010110110001;
            15'd27129: log10_cal = 16'b0000010110110001;
            15'd27130: log10_cal = 16'b0000010110110001;
            15'd27131: log10_cal = 16'b0000010110110001;
            15'd27132: log10_cal = 16'b0000010110110001;
            15'd27133: log10_cal = 16'b0000010110110001;
            15'd27134: log10_cal = 16'b0000010110110001;
            15'd27135: log10_cal = 16'b0000010110110001;
            15'd27136: log10_cal = 16'b0000010110110001;
            15'd27137: log10_cal = 16'b0000010110110001;
            15'd27138: log10_cal = 16'b0000010110110001;
            15'd27139: log10_cal = 16'b0000010110110001;
            15'd27140: log10_cal = 16'b0000010110110001;
            15'd27141: log10_cal = 16'b0000010110110001;
            15'd27142: log10_cal = 16'b0000010110110001;
            15'd27143: log10_cal = 16'b0000010110110001;
            15'd27144: log10_cal = 16'b0000010110110001;
            15'd27145: log10_cal = 16'b0000010110110001;
            15'd27146: log10_cal = 16'b0000010110110001;
            15'd27147: log10_cal = 16'b0000010110110001;
            15'd27148: log10_cal = 16'b0000010110110001;
            15'd27149: log10_cal = 16'b0000010110110001;
            15'd27150: log10_cal = 16'b0000010110110001;
            15'd27151: log10_cal = 16'b0000010110110001;
            15'd27152: log10_cal = 16'b0000010110110001;
            15'd27153: log10_cal = 16'b0000010110110001;
            15'd27154: log10_cal = 16'b0000010110110001;
            15'd27155: log10_cal = 16'b0000010110110001;
            15'd27156: log10_cal = 16'b0000010110110001;
            15'd27157: log10_cal = 16'b0000010110110001;
            15'd27158: log10_cal = 16'b0000010110110001;
            15'd27159: log10_cal = 16'b0000010110110001;
            15'd27160: log10_cal = 16'b0000010110110001;
            15'd27161: log10_cal = 16'b0000010110110001;
            15'd27162: log10_cal = 16'b0000010110110001;
            15'd27163: log10_cal = 16'b0000010110110001;
            15'd27164: log10_cal = 16'b0000010110110001;
            15'd27165: log10_cal = 16'b0000010110110001;
            15'd27166: log10_cal = 16'b0000010110110001;
            15'd27167: log10_cal = 16'b0000010110110001;
            15'd27168: log10_cal = 16'b0000010110110001;
            15'd27169: log10_cal = 16'b0000010110110001;
            15'd27170: log10_cal = 16'b0000010110110001;
            15'd27171: log10_cal = 16'b0000010110110001;
            15'd27172: log10_cal = 16'b0000010110110001;
            15'd27173: log10_cal = 16'b0000010110110010;
            15'd27174: log10_cal = 16'b0000010110110010;
            15'd27175: log10_cal = 16'b0000010110110010;
            15'd27176: log10_cal = 16'b0000010110110010;
            15'd27177: log10_cal = 16'b0000010110110010;
            15'd27178: log10_cal = 16'b0000010110110010;
            15'd27179: log10_cal = 16'b0000010110110010;
            15'd27180: log10_cal = 16'b0000010110110010;
            15'd27181: log10_cal = 16'b0000010110110010;
            15'd27182: log10_cal = 16'b0000010110110010;
            15'd27183: log10_cal = 16'b0000010110110010;
            15'd27184: log10_cal = 16'b0000010110110010;
            15'd27185: log10_cal = 16'b0000010110110010;
            15'd27186: log10_cal = 16'b0000010110110010;
            15'd27187: log10_cal = 16'b0000010110110010;
            15'd27188: log10_cal = 16'b0000010110110010;
            15'd27189: log10_cal = 16'b0000010110110010;
            15'd27190: log10_cal = 16'b0000010110110010;
            15'd27191: log10_cal = 16'b0000010110110010;
            15'd27192: log10_cal = 16'b0000010110110010;
            15'd27193: log10_cal = 16'b0000010110110010;
            15'd27194: log10_cal = 16'b0000010110110010;
            15'd27195: log10_cal = 16'b0000010110110010;
            15'd27196: log10_cal = 16'b0000010110110010;
            15'd27197: log10_cal = 16'b0000010110110010;
            15'd27198: log10_cal = 16'b0000010110110010;
            15'd27199: log10_cal = 16'b0000010110110010;
            15'd27200: log10_cal = 16'b0000010110110010;
            15'd27201: log10_cal = 16'b0000010110110010;
            15'd27202: log10_cal = 16'b0000010110110010;
            15'd27203: log10_cal = 16'b0000010110110010;
            15'd27204: log10_cal = 16'b0000010110110010;
            15'd27205: log10_cal = 16'b0000010110110010;
            15'd27206: log10_cal = 16'b0000010110110010;
            15'd27207: log10_cal = 16'b0000010110110010;
            15'd27208: log10_cal = 16'b0000010110110010;
            15'd27209: log10_cal = 16'b0000010110110010;
            15'd27210: log10_cal = 16'b0000010110110010;
            15'd27211: log10_cal = 16'b0000010110110010;
            15'd27212: log10_cal = 16'b0000010110110010;
            15'd27213: log10_cal = 16'b0000010110110010;
            15'd27214: log10_cal = 16'b0000010110110010;
            15'd27215: log10_cal = 16'b0000010110110010;
            15'd27216: log10_cal = 16'b0000010110110010;
            15'd27217: log10_cal = 16'b0000010110110010;
            15'd27218: log10_cal = 16'b0000010110110010;
            15'd27219: log10_cal = 16'b0000010110110010;
            15'd27220: log10_cal = 16'b0000010110110010;
            15'd27221: log10_cal = 16'b0000010110110010;
            15'd27222: log10_cal = 16'b0000010110110010;
            15'd27223: log10_cal = 16'b0000010110110010;
            15'd27224: log10_cal = 16'b0000010110110010;
            15'd27225: log10_cal = 16'b0000010110110010;
            15'd27226: log10_cal = 16'b0000010110110010;
            15'd27227: log10_cal = 16'b0000010110110010;
            15'd27228: log10_cal = 16'b0000010110110010;
            15'd27229: log10_cal = 16'b0000010110110010;
            15'd27230: log10_cal = 16'b0000010110110010;
            15'd27231: log10_cal = 16'b0000010110110010;
            15'd27232: log10_cal = 16'b0000010110110010;
            15'd27233: log10_cal = 16'b0000010110110010;
            15'd27234: log10_cal = 16'b0000010110110011;
            15'd27235: log10_cal = 16'b0000010110110011;
            15'd27236: log10_cal = 16'b0000010110110011;
            15'd27237: log10_cal = 16'b0000010110110011;
            15'd27238: log10_cal = 16'b0000010110110011;
            15'd27239: log10_cal = 16'b0000010110110011;
            15'd27240: log10_cal = 16'b0000010110110011;
            15'd27241: log10_cal = 16'b0000010110110011;
            15'd27242: log10_cal = 16'b0000010110110011;
            15'd27243: log10_cal = 16'b0000010110110011;
            15'd27244: log10_cal = 16'b0000010110110011;
            15'd27245: log10_cal = 16'b0000010110110011;
            15'd27246: log10_cal = 16'b0000010110110011;
            15'd27247: log10_cal = 16'b0000010110110011;
            15'd27248: log10_cal = 16'b0000010110110011;
            15'd27249: log10_cal = 16'b0000010110110011;
            15'd27250: log10_cal = 16'b0000010110110011;
            15'd27251: log10_cal = 16'b0000010110110011;
            15'd27252: log10_cal = 16'b0000010110110011;
            15'd27253: log10_cal = 16'b0000010110110011;
            15'd27254: log10_cal = 16'b0000010110110011;
            15'd27255: log10_cal = 16'b0000010110110011;
            15'd27256: log10_cal = 16'b0000010110110011;
            15'd27257: log10_cal = 16'b0000010110110011;
            15'd27258: log10_cal = 16'b0000010110110011;
            15'd27259: log10_cal = 16'b0000010110110011;
            15'd27260: log10_cal = 16'b0000010110110011;
            15'd27261: log10_cal = 16'b0000010110110011;
            15'd27262: log10_cal = 16'b0000010110110011;
            15'd27263: log10_cal = 16'b0000010110110011;
            15'd27264: log10_cal = 16'b0000010110110011;
            15'd27265: log10_cal = 16'b0000010110110011;
            15'd27266: log10_cal = 16'b0000010110110011;
            15'd27267: log10_cal = 16'b0000010110110011;
            15'd27268: log10_cal = 16'b0000010110110011;
            15'd27269: log10_cal = 16'b0000010110110011;
            15'd27270: log10_cal = 16'b0000010110110011;
            15'd27271: log10_cal = 16'b0000010110110011;
            15'd27272: log10_cal = 16'b0000010110110011;
            15'd27273: log10_cal = 16'b0000010110110011;
            15'd27274: log10_cal = 16'b0000010110110011;
            15'd27275: log10_cal = 16'b0000010110110011;
            15'd27276: log10_cal = 16'b0000010110110011;
            15'd27277: log10_cal = 16'b0000010110110011;
            15'd27278: log10_cal = 16'b0000010110110011;
            15'd27279: log10_cal = 16'b0000010110110011;
            15'd27280: log10_cal = 16'b0000010110110011;
            15'd27281: log10_cal = 16'b0000010110110011;
            15'd27282: log10_cal = 16'b0000010110110011;
            15'd27283: log10_cal = 16'b0000010110110011;
            15'd27284: log10_cal = 16'b0000010110110011;
            15'd27285: log10_cal = 16'b0000010110110011;
            15'd27286: log10_cal = 16'b0000010110110011;
            15'd27287: log10_cal = 16'b0000010110110011;
            15'd27288: log10_cal = 16'b0000010110110011;
            15'd27289: log10_cal = 16'b0000010110110011;
            15'd27290: log10_cal = 16'b0000010110110011;
            15'd27291: log10_cal = 16'b0000010110110011;
            15'd27292: log10_cal = 16'b0000010110110011;
            15'd27293: log10_cal = 16'b0000010110110011;
            15'd27294: log10_cal = 16'b0000010110110011;
            15'd27295: log10_cal = 16'b0000010110110100;
            15'd27296: log10_cal = 16'b0000010110110100;
            15'd27297: log10_cal = 16'b0000010110110100;
            15'd27298: log10_cal = 16'b0000010110110100;
            15'd27299: log10_cal = 16'b0000010110110100;
            15'd27300: log10_cal = 16'b0000010110110100;
            15'd27301: log10_cal = 16'b0000010110110100;
            15'd27302: log10_cal = 16'b0000010110110100;
            15'd27303: log10_cal = 16'b0000010110110100;
            15'd27304: log10_cal = 16'b0000010110110100;
            15'd27305: log10_cal = 16'b0000010110110100;
            15'd27306: log10_cal = 16'b0000010110110100;
            15'd27307: log10_cal = 16'b0000010110110100;
            15'd27308: log10_cal = 16'b0000010110110100;
            15'd27309: log10_cal = 16'b0000010110110100;
            15'd27310: log10_cal = 16'b0000010110110100;
            15'd27311: log10_cal = 16'b0000010110110100;
            15'd27312: log10_cal = 16'b0000010110110100;
            15'd27313: log10_cal = 16'b0000010110110100;
            15'd27314: log10_cal = 16'b0000010110110100;
            15'd27315: log10_cal = 16'b0000010110110100;
            15'd27316: log10_cal = 16'b0000010110110100;
            15'd27317: log10_cal = 16'b0000010110110100;
            15'd27318: log10_cal = 16'b0000010110110100;
            15'd27319: log10_cal = 16'b0000010110110100;
            15'd27320: log10_cal = 16'b0000010110110100;
            15'd27321: log10_cal = 16'b0000010110110100;
            15'd27322: log10_cal = 16'b0000010110110100;
            15'd27323: log10_cal = 16'b0000010110110100;
            15'd27324: log10_cal = 16'b0000010110110100;
            15'd27325: log10_cal = 16'b0000010110110100;
            15'd27326: log10_cal = 16'b0000010110110100;
            15'd27327: log10_cal = 16'b0000010110110100;
            15'd27328: log10_cal = 16'b0000010110110100;
            15'd27329: log10_cal = 16'b0000010110110100;
            15'd27330: log10_cal = 16'b0000010110110100;
            15'd27331: log10_cal = 16'b0000010110110100;
            15'd27332: log10_cal = 16'b0000010110110100;
            15'd27333: log10_cal = 16'b0000010110110100;
            15'd27334: log10_cal = 16'b0000010110110100;
            15'd27335: log10_cal = 16'b0000010110110100;
            15'd27336: log10_cal = 16'b0000010110110100;
            15'd27337: log10_cal = 16'b0000010110110100;
            15'd27338: log10_cal = 16'b0000010110110100;
            15'd27339: log10_cal = 16'b0000010110110100;
            15'd27340: log10_cal = 16'b0000010110110100;
            15'd27341: log10_cal = 16'b0000010110110100;
            15'd27342: log10_cal = 16'b0000010110110100;
            15'd27343: log10_cal = 16'b0000010110110100;
            15'd27344: log10_cal = 16'b0000010110110100;
            15'd27345: log10_cal = 16'b0000010110110100;
            15'd27346: log10_cal = 16'b0000010110110100;
            15'd27347: log10_cal = 16'b0000010110110100;
            15'd27348: log10_cal = 16'b0000010110110100;
            15'd27349: log10_cal = 16'b0000010110110100;
            15'd27350: log10_cal = 16'b0000010110110100;
            15'd27351: log10_cal = 16'b0000010110110100;
            15'd27352: log10_cal = 16'b0000010110110100;
            15'd27353: log10_cal = 16'b0000010110110100;
            15'd27354: log10_cal = 16'b0000010110110100;
            15'd27355: log10_cal = 16'b0000010110110100;
            15'd27356: log10_cal = 16'b0000010110110100;
            15'd27357: log10_cal = 16'b0000010110110101;
            15'd27358: log10_cal = 16'b0000010110110101;
            15'd27359: log10_cal = 16'b0000010110110101;
            15'd27360: log10_cal = 16'b0000010110110101;
            15'd27361: log10_cal = 16'b0000010110110101;
            15'd27362: log10_cal = 16'b0000010110110101;
            15'd27363: log10_cal = 16'b0000010110110101;
            15'd27364: log10_cal = 16'b0000010110110101;
            15'd27365: log10_cal = 16'b0000010110110101;
            15'd27366: log10_cal = 16'b0000010110110101;
            15'd27367: log10_cal = 16'b0000010110110101;
            15'd27368: log10_cal = 16'b0000010110110101;
            15'd27369: log10_cal = 16'b0000010110110101;
            15'd27370: log10_cal = 16'b0000010110110101;
            15'd27371: log10_cal = 16'b0000010110110101;
            15'd27372: log10_cal = 16'b0000010110110101;
            15'd27373: log10_cal = 16'b0000010110110101;
            15'd27374: log10_cal = 16'b0000010110110101;
            15'd27375: log10_cal = 16'b0000010110110101;
            15'd27376: log10_cal = 16'b0000010110110101;
            15'd27377: log10_cal = 16'b0000010110110101;
            15'd27378: log10_cal = 16'b0000010110110101;
            15'd27379: log10_cal = 16'b0000010110110101;
            15'd27380: log10_cal = 16'b0000010110110101;
            15'd27381: log10_cal = 16'b0000010110110101;
            15'd27382: log10_cal = 16'b0000010110110101;
            15'd27383: log10_cal = 16'b0000010110110101;
            15'd27384: log10_cal = 16'b0000010110110101;
            15'd27385: log10_cal = 16'b0000010110110101;
            15'd27386: log10_cal = 16'b0000010110110101;
            15'd27387: log10_cal = 16'b0000010110110101;
            15'd27388: log10_cal = 16'b0000010110110101;
            15'd27389: log10_cal = 16'b0000010110110101;
            15'd27390: log10_cal = 16'b0000010110110101;
            15'd27391: log10_cal = 16'b0000010110110101;
            15'd27392: log10_cal = 16'b0000010110110101;
            15'd27393: log10_cal = 16'b0000010110110101;
            15'd27394: log10_cal = 16'b0000010110110101;
            15'd27395: log10_cal = 16'b0000010110110101;
            15'd27396: log10_cal = 16'b0000010110110101;
            15'd27397: log10_cal = 16'b0000010110110101;
            15'd27398: log10_cal = 16'b0000010110110101;
            15'd27399: log10_cal = 16'b0000010110110101;
            15'd27400: log10_cal = 16'b0000010110110101;
            15'd27401: log10_cal = 16'b0000010110110101;
            15'd27402: log10_cal = 16'b0000010110110101;
            15'd27403: log10_cal = 16'b0000010110110101;
            15'd27404: log10_cal = 16'b0000010110110101;
            15'd27405: log10_cal = 16'b0000010110110101;
            15'd27406: log10_cal = 16'b0000010110110101;
            15'd27407: log10_cal = 16'b0000010110110101;
            15'd27408: log10_cal = 16'b0000010110110101;
            15'd27409: log10_cal = 16'b0000010110110101;
            15'd27410: log10_cal = 16'b0000010110110101;
            15'd27411: log10_cal = 16'b0000010110110101;
            15'd27412: log10_cal = 16'b0000010110110101;
            15'd27413: log10_cal = 16'b0000010110110101;
            15'd27414: log10_cal = 16'b0000010110110101;
            15'd27415: log10_cal = 16'b0000010110110101;
            15'd27416: log10_cal = 16'b0000010110110101;
            15'd27417: log10_cal = 16'b0000010110110101;
            15'd27418: log10_cal = 16'b0000010110110110;
            15'd27419: log10_cal = 16'b0000010110110110;
            15'd27420: log10_cal = 16'b0000010110110110;
            15'd27421: log10_cal = 16'b0000010110110110;
            15'd27422: log10_cal = 16'b0000010110110110;
            15'd27423: log10_cal = 16'b0000010110110110;
            15'd27424: log10_cal = 16'b0000010110110110;
            15'd27425: log10_cal = 16'b0000010110110110;
            15'd27426: log10_cal = 16'b0000010110110110;
            15'd27427: log10_cal = 16'b0000010110110110;
            15'd27428: log10_cal = 16'b0000010110110110;
            15'd27429: log10_cal = 16'b0000010110110110;
            15'd27430: log10_cal = 16'b0000010110110110;
            15'd27431: log10_cal = 16'b0000010110110110;
            15'd27432: log10_cal = 16'b0000010110110110;
            15'd27433: log10_cal = 16'b0000010110110110;
            15'd27434: log10_cal = 16'b0000010110110110;
            15'd27435: log10_cal = 16'b0000010110110110;
            15'd27436: log10_cal = 16'b0000010110110110;
            15'd27437: log10_cal = 16'b0000010110110110;
            15'd27438: log10_cal = 16'b0000010110110110;
            15'd27439: log10_cal = 16'b0000010110110110;
            15'd27440: log10_cal = 16'b0000010110110110;
            15'd27441: log10_cal = 16'b0000010110110110;
            15'd27442: log10_cal = 16'b0000010110110110;
            15'd27443: log10_cal = 16'b0000010110110110;
            15'd27444: log10_cal = 16'b0000010110110110;
            15'd27445: log10_cal = 16'b0000010110110110;
            15'd27446: log10_cal = 16'b0000010110110110;
            15'd27447: log10_cal = 16'b0000010110110110;
            15'd27448: log10_cal = 16'b0000010110110110;
            15'd27449: log10_cal = 16'b0000010110110110;
            15'd27450: log10_cal = 16'b0000010110110110;
            15'd27451: log10_cal = 16'b0000010110110110;
            15'd27452: log10_cal = 16'b0000010110110110;
            15'd27453: log10_cal = 16'b0000010110110110;
            15'd27454: log10_cal = 16'b0000010110110110;
            15'd27455: log10_cal = 16'b0000010110110110;
            15'd27456: log10_cal = 16'b0000010110110110;
            15'd27457: log10_cal = 16'b0000010110110110;
            15'd27458: log10_cal = 16'b0000010110110110;
            15'd27459: log10_cal = 16'b0000010110110110;
            15'd27460: log10_cal = 16'b0000010110110110;
            15'd27461: log10_cal = 16'b0000010110110110;
            15'd27462: log10_cal = 16'b0000010110110110;
            15'd27463: log10_cal = 16'b0000010110110110;
            15'd27464: log10_cal = 16'b0000010110110110;
            15'd27465: log10_cal = 16'b0000010110110110;
            15'd27466: log10_cal = 16'b0000010110110110;
            15'd27467: log10_cal = 16'b0000010110110110;
            15'd27468: log10_cal = 16'b0000010110110110;
            15'd27469: log10_cal = 16'b0000010110110110;
            15'd27470: log10_cal = 16'b0000010110110110;
            15'd27471: log10_cal = 16'b0000010110110110;
            15'd27472: log10_cal = 16'b0000010110110110;
            15'd27473: log10_cal = 16'b0000010110110110;
            15'd27474: log10_cal = 16'b0000010110110110;
            15'd27475: log10_cal = 16'b0000010110110110;
            15'd27476: log10_cal = 16'b0000010110110110;
            15'd27477: log10_cal = 16'b0000010110110110;
            15'd27478: log10_cal = 16'b0000010110110110;
            15'd27479: log10_cal = 16'b0000010110110110;
            15'd27480: log10_cal = 16'b0000010110110111;
            15'd27481: log10_cal = 16'b0000010110110111;
            15'd27482: log10_cal = 16'b0000010110110111;
            15'd27483: log10_cal = 16'b0000010110110111;
            15'd27484: log10_cal = 16'b0000010110110111;
            15'd27485: log10_cal = 16'b0000010110110111;
            15'd27486: log10_cal = 16'b0000010110110111;
            15'd27487: log10_cal = 16'b0000010110110111;
            15'd27488: log10_cal = 16'b0000010110110111;
            15'd27489: log10_cal = 16'b0000010110110111;
            15'd27490: log10_cal = 16'b0000010110110111;
            15'd27491: log10_cal = 16'b0000010110110111;
            15'd27492: log10_cal = 16'b0000010110110111;
            15'd27493: log10_cal = 16'b0000010110110111;
            15'd27494: log10_cal = 16'b0000010110110111;
            15'd27495: log10_cal = 16'b0000010110110111;
            15'd27496: log10_cal = 16'b0000010110110111;
            15'd27497: log10_cal = 16'b0000010110110111;
            15'd27498: log10_cal = 16'b0000010110110111;
            15'd27499: log10_cal = 16'b0000010110110111;
            15'd27500: log10_cal = 16'b0000010110110111;
            15'd27501: log10_cal = 16'b0000010110110111;
            15'd27502: log10_cal = 16'b0000010110110111;
            15'd27503: log10_cal = 16'b0000010110110111;
            15'd27504: log10_cal = 16'b0000010110110111;
            15'd27505: log10_cal = 16'b0000010110110111;
            15'd27506: log10_cal = 16'b0000010110110111;
            15'd27507: log10_cal = 16'b0000010110110111;
            15'd27508: log10_cal = 16'b0000010110110111;
            15'd27509: log10_cal = 16'b0000010110110111;
            15'd27510: log10_cal = 16'b0000010110110111;
            15'd27511: log10_cal = 16'b0000010110110111;
            15'd27512: log10_cal = 16'b0000010110110111;
            15'd27513: log10_cal = 16'b0000010110110111;
            15'd27514: log10_cal = 16'b0000010110110111;
            15'd27515: log10_cal = 16'b0000010110110111;
            15'd27516: log10_cal = 16'b0000010110110111;
            15'd27517: log10_cal = 16'b0000010110110111;
            15'd27518: log10_cal = 16'b0000010110110111;
            15'd27519: log10_cal = 16'b0000010110110111;
            15'd27520: log10_cal = 16'b0000010110110111;
            15'd27521: log10_cal = 16'b0000010110110111;
            15'd27522: log10_cal = 16'b0000010110110111;
            15'd27523: log10_cal = 16'b0000010110110111;
            15'd27524: log10_cal = 16'b0000010110110111;
            15'd27525: log10_cal = 16'b0000010110110111;
            15'd27526: log10_cal = 16'b0000010110110111;
            15'd27527: log10_cal = 16'b0000010110110111;
            15'd27528: log10_cal = 16'b0000010110110111;
            15'd27529: log10_cal = 16'b0000010110110111;
            15'd27530: log10_cal = 16'b0000010110110111;
            15'd27531: log10_cal = 16'b0000010110110111;
            15'd27532: log10_cal = 16'b0000010110110111;
            15'd27533: log10_cal = 16'b0000010110110111;
            15'd27534: log10_cal = 16'b0000010110110111;
            15'd27535: log10_cal = 16'b0000010110110111;
            15'd27536: log10_cal = 16'b0000010110110111;
            15'd27537: log10_cal = 16'b0000010110110111;
            15'd27538: log10_cal = 16'b0000010110110111;
            15'd27539: log10_cal = 16'b0000010110110111;
            15'd27540: log10_cal = 16'b0000010110110111;
            15'd27541: log10_cal = 16'b0000010110110111;
            15'd27542: log10_cal = 16'b0000010110111000;
            15'd27543: log10_cal = 16'b0000010110111000;
            15'd27544: log10_cal = 16'b0000010110111000;
            15'd27545: log10_cal = 16'b0000010110111000;
            15'd27546: log10_cal = 16'b0000010110111000;
            15'd27547: log10_cal = 16'b0000010110111000;
            15'd27548: log10_cal = 16'b0000010110111000;
            15'd27549: log10_cal = 16'b0000010110111000;
            15'd27550: log10_cal = 16'b0000010110111000;
            15'd27551: log10_cal = 16'b0000010110111000;
            15'd27552: log10_cal = 16'b0000010110111000;
            15'd27553: log10_cal = 16'b0000010110111000;
            15'd27554: log10_cal = 16'b0000010110111000;
            15'd27555: log10_cal = 16'b0000010110111000;
            15'd27556: log10_cal = 16'b0000010110111000;
            15'd27557: log10_cal = 16'b0000010110111000;
            15'd27558: log10_cal = 16'b0000010110111000;
            15'd27559: log10_cal = 16'b0000010110111000;
            15'd27560: log10_cal = 16'b0000010110111000;
            15'd27561: log10_cal = 16'b0000010110111000;
            15'd27562: log10_cal = 16'b0000010110111000;
            15'd27563: log10_cal = 16'b0000010110111000;
            15'd27564: log10_cal = 16'b0000010110111000;
            15'd27565: log10_cal = 16'b0000010110111000;
            15'd27566: log10_cal = 16'b0000010110111000;
            15'd27567: log10_cal = 16'b0000010110111000;
            15'd27568: log10_cal = 16'b0000010110111000;
            15'd27569: log10_cal = 16'b0000010110111000;
            15'd27570: log10_cal = 16'b0000010110111000;
            15'd27571: log10_cal = 16'b0000010110111000;
            15'd27572: log10_cal = 16'b0000010110111000;
            15'd27573: log10_cal = 16'b0000010110111000;
            15'd27574: log10_cal = 16'b0000010110111000;
            15'd27575: log10_cal = 16'b0000010110111000;
            15'd27576: log10_cal = 16'b0000010110111000;
            15'd27577: log10_cal = 16'b0000010110111000;
            15'd27578: log10_cal = 16'b0000010110111000;
            15'd27579: log10_cal = 16'b0000010110111000;
            15'd27580: log10_cal = 16'b0000010110111000;
            15'd27581: log10_cal = 16'b0000010110111000;
            15'd27582: log10_cal = 16'b0000010110111000;
            15'd27583: log10_cal = 16'b0000010110111000;
            15'd27584: log10_cal = 16'b0000010110111000;
            15'd27585: log10_cal = 16'b0000010110111000;
            15'd27586: log10_cal = 16'b0000010110111000;
            15'd27587: log10_cal = 16'b0000010110111000;
            15'd27588: log10_cal = 16'b0000010110111000;
            15'd27589: log10_cal = 16'b0000010110111000;
            15'd27590: log10_cal = 16'b0000010110111000;
            15'd27591: log10_cal = 16'b0000010110111000;
            15'd27592: log10_cal = 16'b0000010110111000;
            15'd27593: log10_cal = 16'b0000010110111000;
            15'd27594: log10_cal = 16'b0000010110111000;
            15'd27595: log10_cal = 16'b0000010110111000;
            15'd27596: log10_cal = 16'b0000010110111000;
            15'd27597: log10_cal = 16'b0000010110111000;
            15'd27598: log10_cal = 16'b0000010110111000;
            15'd27599: log10_cal = 16'b0000010110111000;
            15'd27600: log10_cal = 16'b0000010110111000;
            15'd27601: log10_cal = 16'b0000010110111000;
            15'd27602: log10_cal = 16'b0000010110111000;
            15'd27603: log10_cal = 16'b0000010110111000;
            15'd27604: log10_cal = 16'b0000010110111001;
            15'd27605: log10_cal = 16'b0000010110111001;
            15'd27606: log10_cal = 16'b0000010110111001;
            15'd27607: log10_cal = 16'b0000010110111001;
            15'd27608: log10_cal = 16'b0000010110111001;
            15'd27609: log10_cal = 16'b0000010110111001;
            15'd27610: log10_cal = 16'b0000010110111001;
            15'd27611: log10_cal = 16'b0000010110111001;
            15'd27612: log10_cal = 16'b0000010110111001;
            15'd27613: log10_cal = 16'b0000010110111001;
            15'd27614: log10_cal = 16'b0000010110111001;
            15'd27615: log10_cal = 16'b0000010110111001;
            15'd27616: log10_cal = 16'b0000010110111001;
            15'd27617: log10_cal = 16'b0000010110111001;
            15'd27618: log10_cal = 16'b0000010110111001;
            15'd27619: log10_cal = 16'b0000010110111001;
            15'd27620: log10_cal = 16'b0000010110111001;
            15'd27621: log10_cal = 16'b0000010110111001;
            15'd27622: log10_cal = 16'b0000010110111001;
            15'd27623: log10_cal = 16'b0000010110111001;
            15'd27624: log10_cal = 16'b0000010110111001;
            15'd27625: log10_cal = 16'b0000010110111001;
            15'd27626: log10_cal = 16'b0000010110111001;
            15'd27627: log10_cal = 16'b0000010110111001;
            15'd27628: log10_cal = 16'b0000010110111001;
            15'd27629: log10_cal = 16'b0000010110111001;
            15'd27630: log10_cal = 16'b0000010110111001;
            15'd27631: log10_cal = 16'b0000010110111001;
            15'd27632: log10_cal = 16'b0000010110111001;
            15'd27633: log10_cal = 16'b0000010110111001;
            15'd27634: log10_cal = 16'b0000010110111001;
            15'd27635: log10_cal = 16'b0000010110111001;
            15'd27636: log10_cal = 16'b0000010110111001;
            15'd27637: log10_cal = 16'b0000010110111001;
            15'd27638: log10_cal = 16'b0000010110111001;
            15'd27639: log10_cal = 16'b0000010110111001;
            15'd27640: log10_cal = 16'b0000010110111001;
            15'd27641: log10_cal = 16'b0000010110111001;
            15'd27642: log10_cal = 16'b0000010110111001;
            15'd27643: log10_cal = 16'b0000010110111001;
            15'd27644: log10_cal = 16'b0000010110111001;
            15'd27645: log10_cal = 16'b0000010110111001;
            15'd27646: log10_cal = 16'b0000010110111001;
            15'd27647: log10_cal = 16'b0000010110111001;
            15'd27648: log10_cal = 16'b0000010110111001;
            15'd27649: log10_cal = 16'b0000010110111001;
            15'd27650: log10_cal = 16'b0000010110111001;
            15'd27651: log10_cal = 16'b0000010110111001;
            15'd27652: log10_cal = 16'b0000010110111001;
            15'd27653: log10_cal = 16'b0000010110111001;
            15'd27654: log10_cal = 16'b0000010110111001;
            15'd27655: log10_cal = 16'b0000010110111001;
            15'd27656: log10_cal = 16'b0000010110111001;
            15'd27657: log10_cal = 16'b0000010110111001;
            15'd27658: log10_cal = 16'b0000010110111001;
            15'd27659: log10_cal = 16'b0000010110111001;
            15'd27660: log10_cal = 16'b0000010110111001;
            15'd27661: log10_cal = 16'b0000010110111001;
            15'd27662: log10_cal = 16'b0000010110111001;
            15'd27663: log10_cal = 16'b0000010110111001;
            15'd27664: log10_cal = 16'b0000010110111001;
            15'd27665: log10_cal = 16'b0000010110111001;
            15'd27666: log10_cal = 16'b0000010110111010;
            15'd27667: log10_cal = 16'b0000010110111010;
            15'd27668: log10_cal = 16'b0000010110111010;
            15'd27669: log10_cal = 16'b0000010110111010;
            15'd27670: log10_cal = 16'b0000010110111010;
            15'd27671: log10_cal = 16'b0000010110111010;
            15'd27672: log10_cal = 16'b0000010110111010;
            15'd27673: log10_cal = 16'b0000010110111010;
            15'd27674: log10_cal = 16'b0000010110111010;
            15'd27675: log10_cal = 16'b0000010110111010;
            15'd27676: log10_cal = 16'b0000010110111010;
            15'd27677: log10_cal = 16'b0000010110111010;
            15'd27678: log10_cal = 16'b0000010110111010;
            15'd27679: log10_cal = 16'b0000010110111010;
            15'd27680: log10_cal = 16'b0000010110111010;
            15'd27681: log10_cal = 16'b0000010110111010;
            15'd27682: log10_cal = 16'b0000010110111010;
            15'd27683: log10_cal = 16'b0000010110111010;
            15'd27684: log10_cal = 16'b0000010110111010;
            15'd27685: log10_cal = 16'b0000010110111010;
            15'd27686: log10_cal = 16'b0000010110111010;
            15'd27687: log10_cal = 16'b0000010110111010;
            15'd27688: log10_cal = 16'b0000010110111010;
            15'd27689: log10_cal = 16'b0000010110111010;
            15'd27690: log10_cal = 16'b0000010110111010;
            15'd27691: log10_cal = 16'b0000010110111010;
            15'd27692: log10_cal = 16'b0000010110111010;
            15'd27693: log10_cal = 16'b0000010110111010;
            15'd27694: log10_cal = 16'b0000010110111010;
            15'd27695: log10_cal = 16'b0000010110111010;
            15'd27696: log10_cal = 16'b0000010110111010;
            15'd27697: log10_cal = 16'b0000010110111010;
            15'd27698: log10_cal = 16'b0000010110111010;
            15'd27699: log10_cal = 16'b0000010110111010;
            15'd27700: log10_cal = 16'b0000010110111010;
            15'd27701: log10_cal = 16'b0000010110111010;
            15'd27702: log10_cal = 16'b0000010110111010;
            15'd27703: log10_cal = 16'b0000010110111010;
            15'd27704: log10_cal = 16'b0000010110111010;
            15'd27705: log10_cal = 16'b0000010110111010;
            15'd27706: log10_cal = 16'b0000010110111010;
            15'd27707: log10_cal = 16'b0000010110111010;
            15'd27708: log10_cal = 16'b0000010110111010;
            15'd27709: log10_cal = 16'b0000010110111010;
            15'd27710: log10_cal = 16'b0000010110111010;
            15'd27711: log10_cal = 16'b0000010110111010;
            15'd27712: log10_cal = 16'b0000010110111010;
            15'd27713: log10_cal = 16'b0000010110111010;
            15'd27714: log10_cal = 16'b0000010110111010;
            15'd27715: log10_cal = 16'b0000010110111010;
            15'd27716: log10_cal = 16'b0000010110111010;
            15'd27717: log10_cal = 16'b0000010110111010;
            15'd27718: log10_cal = 16'b0000010110111010;
            15'd27719: log10_cal = 16'b0000010110111010;
            15'd27720: log10_cal = 16'b0000010110111010;
            15'd27721: log10_cal = 16'b0000010110111010;
            15'd27722: log10_cal = 16'b0000010110111010;
            15'd27723: log10_cal = 16'b0000010110111010;
            15'd27724: log10_cal = 16'b0000010110111010;
            15'd27725: log10_cal = 16'b0000010110111010;
            15'd27726: log10_cal = 16'b0000010110111010;
            15'd27727: log10_cal = 16'b0000010110111010;
            15'd27728: log10_cal = 16'b0000010110111011;
            15'd27729: log10_cal = 16'b0000010110111011;
            15'd27730: log10_cal = 16'b0000010110111011;
            15'd27731: log10_cal = 16'b0000010110111011;
            15'd27732: log10_cal = 16'b0000010110111011;
            15'd27733: log10_cal = 16'b0000010110111011;
            15'd27734: log10_cal = 16'b0000010110111011;
            15'd27735: log10_cal = 16'b0000010110111011;
            15'd27736: log10_cal = 16'b0000010110111011;
            15'd27737: log10_cal = 16'b0000010110111011;
            15'd27738: log10_cal = 16'b0000010110111011;
            15'd27739: log10_cal = 16'b0000010110111011;
            15'd27740: log10_cal = 16'b0000010110111011;
            15'd27741: log10_cal = 16'b0000010110111011;
            15'd27742: log10_cal = 16'b0000010110111011;
            15'd27743: log10_cal = 16'b0000010110111011;
            15'd27744: log10_cal = 16'b0000010110111011;
            15'd27745: log10_cal = 16'b0000010110111011;
            15'd27746: log10_cal = 16'b0000010110111011;
            15'd27747: log10_cal = 16'b0000010110111011;
            15'd27748: log10_cal = 16'b0000010110111011;
            15'd27749: log10_cal = 16'b0000010110111011;
            15'd27750: log10_cal = 16'b0000010110111011;
            15'd27751: log10_cal = 16'b0000010110111011;
            15'd27752: log10_cal = 16'b0000010110111011;
            15'd27753: log10_cal = 16'b0000010110111011;
            15'd27754: log10_cal = 16'b0000010110111011;
            15'd27755: log10_cal = 16'b0000010110111011;
            15'd27756: log10_cal = 16'b0000010110111011;
            15'd27757: log10_cal = 16'b0000010110111011;
            15'd27758: log10_cal = 16'b0000010110111011;
            15'd27759: log10_cal = 16'b0000010110111011;
            15'd27760: log10_cal = 16'b0000010110111011;
            15'd27761: log10_cal = 16'b0000010110111011;
            15'd27762: log10_cal = 16'b0000010110111011;
            15'd27763: log10_cal = 16'b0000010110111011;
            15'd27764: log10_cal = 16'b0000010110111011;
            15'd27765: log10_cal = 16'b0000010110111011;
            15'd27766: log10_cal = 16'b0000010110111011;
            15'd27767: log10_cal = 16'b0000010110111011;
            15'd27768: log10_cal = 16'b0000010110111011;
            15'd27769: log10_cal = 16'b0000010110111011;
            15'd27770: log10_cal = 16'b0000010110111011;
            15'd27771: log10_cal = 16'b0000010110111011;
            15'd27772: log10_cal = 16'b0000010110111011;
            15'd27773: log10_cal = 16'b0000010110111011;
            15'd27774: log10_cal = 16'b0000010110111011;
            15'd27775: log10_cal = 16'b0000010110111011;
            15'd27776: log10_cal = 16'b0000010110111011;
            15'd27777: log10_cal = 16'b0000010110111011;
            15'd27778: log10_cal = 16'b0000010110111011;
            15'd27779: log10_cal = 16'b0000010110111011;
            15'd27780: log10_cal = 16'b0000010110111011;
            15'd27781: log10_cal = 16'b0000010110111011;
            15'd27782: log10_cal = 16'b0000010110111011;
            15'd27783: log10_cal = 16'b0000010110111011;
            15'd27784: log10_cal = 16'b0000010110111011;
            15'd27785: log10_cal = 16'b0000010110111011;
            15'd27786: log10_cal = 16'b0000010110111011;
            15'd27787: log10_cal = 16'b0000010110111011;
            15'd27788: log10_cal = 16'b0000010110111011;
            15'd27789: log10_cal = 16'b0000010110111011;
            15'd27790: log10_cal = 16'b0000010110111011;
            15'd27791: log10_cal = 16'b0000010110111100;
            15'd27792: log10_cal = 16'b0000010110111100;
            15'd27793: log10_cal = 16'b0000010110111100;
            15'd27794: log10_cal = 16'b0000010110111100;
            15'd27795: log10_cal = 16'b0000010110111100;
            15'd27796: log10_cal = 16'b0000010110111100;
            15'd27797: log10_cal = 16'b0000010110111100;
            15'd27798: log10_cal = 16'b0000010110111100;
            15'd27799: log10_cal = 16'b0000010110111100;
            15'd27800: log10_cal = 16'b0000010110111100;
            15'd27801: log10_cal = 16'b0000010110111100;
            15'd27802: log10_cal = 16'b0000010110111100;
            15'd27803: log10_cal = 16'b0000010110111100;
            15'd27804: log10_cal = 16'b0000010110111100;
            15'd27805: log10_cal = 16'b0000010110111100;
            15'd27806: log10_cal = 16'b0000010110111100;
            15'd27807: log10_cal = 16'b0000010110111100;
            15'd27808: log10_cal = 16'b0000010110111100;
            15'd27809: log10_cal = 16'b0000010110111100;
            15'd27810: log10_cal = 16'b0000010110111100;
            15'd27811: log10_cal = 16'b0000010110111100;
            15'd27812: log10_cal = 16'b0000010110111100;
            15'd27813: log10_cal = 16'b0000010110111100;
            15'd27814: log10_cal = 16'b0000010110111100;
            15'd27815: log10_cal = 16'b0000010110111100;
            15'd27816: log10_cal = 16'b0000010110111100;
            15'd27817: log10_cal = 16'b0000010110111100;
            15'd27818: log10_cal = 16'b0000010110111100;
            15'd27819: log10_cal = 16'b0000010110111100;
            15'd27820: log10_cal = 16'b0000010110111100;
            15'd27821: log10_cal = 16'b0000010110111100;
            15'd27822: log10_cal = 16'b0000010110111100;
            15'd27823: log10_cal = 16'b0000010110111100;
            15'd27824: log10_cal = 16'b0000010110111100;
            15'd27825: log10_cal = 16'b0000010110111100;
            15'd27826: log10_cal = 16'b0000010110111100;
            15'd27827: log10_cal = 16'b0000010110111100;
            15'd27828: log10_cal = 16'b0000010110111100;
            15'd27829: log10_cal = 16'b0000010110111100;
            15'd27830: log10_cal = 16'b0000010110111100;
            15'd27831: log10_cal = 16'b0000010110111100;
            15'd27832: log10_cal = 16'b0000010110111100;
            15'd27833: log10_cal = 16'b0000010110111100;
            15'd27834: log10_cal = 16'b0000010110111100;
            15'd27835: log10_cal = 16'b0000010110111100;
            15'd27836: log10_cal = 16'b0000010110111100;
            15'd27837: log10_cal = 16'b0000010110111100;
            15'd27838: log10_cal = 16'b0000010110111100;
            15'd27839: log10_cal = 16'b0000010110111100;
            15'd27840: log10_cal = 16'b0000010110111100;
            15'd27841: log10_cal = 16'b0000010110111100;
            15'd27842: log10_cal = 16'b0000010110111100;
            15'd27843: log10_cal = 16'b0000010110111100;
            15'd27844: log10_cal = 16'b0000010110111100;
            15'd27845: log10_cal = 16'b0000010110111100;
            15'd27846: log10_cal = 16'b0000010110111100;
            15'd27847: log10_cal = 16'b0000010110111100;
            15'd27848: log10_cal = 16'b0000010110111100;
            15'd27849: log10_cal = 16'b0000010110111100;
            15'd27850: log10_cal = 16'b0000010110111100;
            15'd27851: log10_cal = 16'b0000010110111100;
            15'd27852: log10_cal = 16'b0000010110111100;
            15'd27853: log10_cal = 16'b0000010110111101;
            15'd27854: log10_cal = 16'b0000010110111101;
            15'd27855: log10_cal = 16'b0000010110111101;
            15'd27856: log10_cal = 16'b0000010110111101;
            15'd27857: log10_cal = 16'b0000010110111101;
            15'd27858: log10_cal = 16'b0000010110111101;
            15'd27859: log10_cal = 16'b0000010110111101;
            15'd27860: log10_cal = 16'b0000010110111101;
            15'd27861: log10_cal = 16'b0000010110111101;
            15'd27862: log10_cal = 16'b0000010110111101;
            15'd27863: log10_cal = 16'b0000010110111101;
            15'd27864: log10_cal = 16'b0000010110111101;
            15'd27865: log10_cal = 16'b0000010110111101;
            15'd27866: log10_cal = 16'b0000010110111101;
            15'd27867: log10_cal = 16'b0000010110111101;
            15'd27868: log10_cal = 16'b0000010110111101;
            15'd27869: log10_cal = 16'b0000010110111101;
            15'd27870: log10_cal = 16'b0000010110111101;
            15'd27871: log10_cal = 16'b0000010110111101;
            15'd27872: log10_cal = 16'b0000010110111101;
            15'd27873: log10_cal = 16'b0000010110111101;
            15'd27874: log10_cal = 16'b0000010110111101;
            15'd27875: log10_cal = 16'b0000010110111101;
            15'd27876: log10_cal = 16'b0000010110111101;
            15'd27877: log10_cal = 16'b0000010110111101;
            15'd27878: log10_cal = 16'b0000010110111101;
            15'd27879: log10_cal = 16'b0000010110111101;
            15'd27880: log10_cal = 16'b0000010110111101;
            15'd27881: log10_cal = 16'b0000010110111101;
            15'd27882: log10_cal = 16'b0000010110111101;
            15'd27883: log10_cal = 16'b0000010110111101;
            15'd27884: log10_cal = 16'b0000010110111101;
            15'd27885: log10_cal = 16'b0000010110111101;
            15'd27886: log10_cal = 16'b0000010110111101;
            15'd27887: log10_cal = 16'b0000010110111101;
            15'd27888: log10_cal = 16'b0000010110111101;
            15'd27889: log10_cal = 16'b0000010110111101;
            15'd27890: log10_cal = 16'b0000010110111101;
            15'd27891: log10_cal = 16'b0000010110111101;
            15'd27892: log10_cal = 16'b0000010110111101;
            15'd27893: log10_cal = 16'b0000010110111101;
            15'd27894: log10_cal = 16'b0000010110111101;
            15'd27895: log10_cal = 16'b0000010110111101;
            15'd27896: log10_cal = 16'b0000010110111101;
            15'd27897: log10_cal = 16'b0000010110111101;
            15'd27898: log10_cal = 16'b0000010110111101;
            15'd27899: log10_cal = 16'b0000010110111101;
            15'd27900: log10_cal = 16'b0000010110111101;
            15'd27901: log10_cal = 16'b0000010110111101;
            15'd27902: log10_cal = 16'b0000010110111101;
            15'd27903: log10_cal = 16'b0000010110111101;
            15'd27904: log10_cal = 16'b0000010110111101;
            15'd27905: log10_cal = 16'b0000010110111101;
            15'd27906: log10_cal = 16'b0000010110111101;
            15'd27907: log10_cal = 16'b0000010110111101;
            15'd27908: log10_cal = 16'b0000010110111101;
            15'd27909: log10_cal = 16'b0000010110111101;
            15'd27910: log10_cal = 16'b0000010110111101;
            15'd27911: log10_cal = 16'b0000010110111101;
            15'd27912: log10_cal = 16'b0000010110111101;
            15'd27913: log10_cal = 16'b0000010110111101;
            15'd27914: log10_cal = 16'b0000010110111101;
            15'd27915: log10_cal = 16'b0000010110111101;
            15'd27916: log10_cal = 16'b0000010110111110;
            15'd27917: log10_cal = 16'b0000010110111110;
            15'd27918: log10_cal = 16'b0000010110111110;
            15'd27919: log10_cal = 16'b0000010110111110;
            15'd27920: log10_cal = 16'b0000010110111110;
            15'd27921: log10_cal = 16'b0000010110111110;
            15'd27922: log10_cal = 16'b0000010110111110;
            15'd27923: log10_cal = 16'b0000010110111110;
            15'd27924: log10_cal = 16'b0000010110111110;
            15'd27925: log10_cal = 16'b0000010110111110;
            15'd27926: log10_cal = 16'b0000010110111110;
            15'd27927: log10_cal = 16'b0000010110111110;
            15'd27928: log10_cal = 16'b0000010110111110;
            15'd27929: log10_cal = 16'b0000010110111110;
            15'd27930: log10_cal = 16'b0000010110111110;
            15'd27931: log10_cal = 16'b0000010110111110;
            15'd27932: log10_cal = 16'b0000010110111110;
            15'd27933: log10_cal = 16'b0000010110111110;
            15'd27934: log10_cal = 16'b0000010110111110;
            15'd27935: log10_cal = 16'b0000010110111110;
            15'd27936: log10_cal = 16'b0000010110111110;
            15'd27937: log10_cal = 16'b0000010110111110;
            15'd27938: log10_cal = 16'b0000010110111110;
            15'd27939: log10_cal = 16'b0000010110111110;
            15'd27940: log10_cal = 16'b0000010110111110;
            15'd27941: log10_cal = 16'b0000010110111110;
            15'd27942: log10_cal = 16'b0000010110111110;
            15'd27943: log10_cal = 16'b0000010110111110;
            15'd27944: log10_cal = 16'b0000010110111110;
            15'd27945: log10_cal = 16'b0000010110111110;
            15'd27946: log10_cal = 16'b0000010110111110;
            15'd27947: log10_cal = 16'b0000010110111110;
            15'd27948: log10_cal = 16'b0000010110111110;
            15'd27949: log10_cal = 16'b0000010110111110;
            15'd27950: log10_cal = 16'b0000010110111110;
            15'd27951: log10_cal = 16'b0000010110111110;
            15'd27952: log10_cal = 16'b0000010110111110;
            15'd27953: log10_cal = 16'b0000010110111110;
            15'd27954: log10_cal = 16'b0000010110111110;
            15'd27955: log10_cal = 16'b0000010110111110;
            15'd27956: log10_cal = 16'b0000010110111110;
            15'd27957: log10_cal = 16'b0000010110111110;
            15'd27958: log10_cal = 16'b0000010110111110;
            15'd27959: log10_cal = 16'b0000010110111110;
            15'd27960: log10_cal = 16'b0000010110111110;
            15'd27961: log10_cal = 16'b0000010110111110;
            15'd27962: log10_cal = 16'b0000010110111110;
            15'd27963: log10_cal = 16'b0000010110111110;
            15'd27964: log10_cal = 16'b0000010110111110;
            15'd27965: log10_cal = 16'b0000010110111110;
            15'd27966: log10_cal = 16'b0000010110111110;
            15'd27967: log10_cal = 16'b0000010110111110;
            15'd27968: log10_cal = 16'b0000010110111110;
            15'd27969: log10_cal = 16'b0000010110111110;
            15'd27970: log10_cal = 16'b0000010110111110;
            15'd27971: log10_cal = 16'b0000010110111110;
            15'd27972: log10_cal = 16'b0000010110111110;
            15'd27973: log10_cal = 16'b0000010110111110;
            15'd27974: log10_cal = 16'b0000010110111110;
            15'd27975: log10_cal = 16'b0000010110111110;
            15'd27976: log10_cal = 16'b0000010110111110;
            15'd27977: log10_cal = 16'b0000010110111110;
            15'd27978: log10_cal = 16'b0000010110111110;
            15'd27979: log10_cal = 16'b0000010110111111;
            15'd27980: log10_cal = 16'b0000010110111111;
            15'd27981: log10_cal = 16'b0000010110111111;
            15'd27982: log10_cal = 16'b0000010110111111;
            15'd27983: log10_cal = 16'b0000010110111111;
            15'd27984: log10_cal = 16'b0000010110111111;
            15'd27985: log10_cal = 16'b0000010110111111;
            15'd27986: log10_cal = 16'b0000010110111111;
            15'd27987: log10_cal = 16'b0000010110111111;
            15'd27988: log10_cal = 16'b0000010110111111;
            15'd27989: log10_cal = 16'b0000010110111111;
            15'd27990: log10_cal = 16'b0000010110111111;
            15'd27991: log10_cal = 16'b0000010110111111;
            15'd27992: log10_cal = 16'b0000010110111111;
            15'd27993: log10_cal = 16'b0000010110111111;
            15'd27994: log10_cal = 16'b0000010110111111;
            15'd27995: log10_cal = 16'b0000010110111111;
            15'd27996: log10_cal = 16'b0000010110111111;
            15'd27997: log10_cal = 16'b0000010110111111;
            15'd27998: log10_cal = 16'b0000010110111111;
            15'd27999: log10_cal = 16'b0000010110111111;
            15'd28000: log10_cal = 16'b0000010110111111;
            15'd28001: log10_cal = 16'b0000010110111111;
            15'd28002: log10_cal = 16'b0000010110111111;
            15'd28003: log10_cal = 16'b0000010110111111;
            15'd28004: log10_cal = 16'b0000010110111111;
            15'd28005: log10_cal = 16'b0000010110111111;
            15'd28006: log10_cal = 16'b0000010110111111;
            15'd28007: log10_cal = 16'b0000010110111111;
            15'd28008: log10_cal = 16'b0000010110111111;
            15'd28009: log10_cal = 16'b0000010110111111;
            15'd28010: log10_cal = 16'b0000010110111111;
            15'd28011: log10_cal = 16'b0000010110111111;
            15'd28012: log10_cal = 16'b0000010110111111;
            15'd28013: log10_cal = 16'b0000010110111111;
            15'd28014: log10_cal = 16'b0000010110111111;
            15'd28015: log10_cal = 16'b0000010110111111;
            15'd28016: log10_cal = 16'b0000010110111111;
            15'd28017: log10_cal = 16'b0000010110111111;
            15'd28018: log10_cal = 16'b0000010110111111;
            15'd28019: log10_cal = 16'b0000010110111111;
            15'd28020: log10_cal = 16'b0000010110111111;
            15'd28021: log10_cal = 16'b0000010110111111;
            15'd28022: log10_cal = 16'b0000010110111111;
            15'd28023: log10_cal = 16'b0000010110111111;
            15'd28024: log10_cal = 16'b0000010110111111;
            15'd28025: log10_cal = 16'b0000010110111111;
            15'd28026: log10_cal = 16'b0000010110111111;
            15'd28027: log10_cal = 16'b0000010110111111;
            15'd28028: log10_cal = 16'b0000010110111111;
            15'd28029: log10_cal = 16'b0000010110111111;
            15'd28030: log10_cal = 16'b0000010110111111;
            15'd28031: log10_cal = 16'b0000010110111111;
            15'd28032: log10_cal = 16'b0000010110111111;
            15'd28033: log10_cal = 16'b0000010110111111;
            15'd28034: log10_cal = 16'b0000010110111111;
            15'd28035: log10_cal = 16'b0000010110111111;
            15'd28036: log10_cal = 16'b0000010110111111;
            15'd28037: log10_cal = 16'b0000010110111111;
            15'd28038: log10_cal = 16'b0000010110111111;
            15'd28039: log10_cal = 16'b0000010110111111;
            15'd28040: log10_cal = 16'b0000010110111111;
            15'd28041: log10_cal = 16'b0000010110111111;
            15'd28042: log10_cal = 16'b0000010111000000;
            15'd28043: log10_cal = 16'b0000010111000000;
            15'd28044: log10_cal = 16'b0000010111000000;
            15'd28045: log10_cal = 16'b0000010111000000;
            15'd28046: log10_cal = 16'b0000010111000000;
            15'd28047: log10_cal = 16'b0000010111000000;
            15'd28048: log10_cal = 16'b0000010111000000;
            15'd28049: log10_cal = 16'b0000010111000000;
            15'd28050: log10_cal = 16'b0000010111000000;
            15'd28051: log10_cal = 16'b0000010111000000;
            15'd28052: log10_cal = 16'b0000010111000000;
            15'd28053: log10_cal = 16'b0000010111000000;
            15'd28054: log10_cal = 16'b0000010111000000;
            15'd28055: log10_cal = 16'b0000010111000000;
            15'd28056: log10_cal = 16'b0000010111000000;
            15'd28057: log10_cal = 16'b0000010111000000;
            15'd28058: log10_cal = 16'b0000010111000000;
            15'd28059: log10_cal = 16'b0000010111000000;
            15'd28060: log10_cal = 16'b0000010111000000;
            15'd28061: log10_cal = 16'b0000010111000000;
            15'd28062: log10_cal = 16'b0000010111000000;
            15'd28063: log10_cal = 16'b0000010111000000;
            15'd28064: log10_cal = 16'b0000010111000000;
            15'd28065: log10_cal = 16'b0000010111000000;
            15'd28066: log10_cal = 16'b0000010111000000;
            15'd28067: log10_cal = 16'b0000010111000000;
            15'd28068: log10_cal = 16'b0000010111000000;
            15'd28069: log10_cal = 16'b0000010111000000;
            15'd28070: log10_cal = 16'b0000010111000000;
            15'd28071: log10_cal = 16'b0000010111000000;
            15'd28072: log10_cal = 16'b0000010111000000;
            15'd28073: log10_cal = 16'b0000010111000000;
            15'd28074: log10_cal = 16'b0000010111000000;
            15'd28075: log10_cal = 16'b0000010111000000;
            15'd28076: log10_cal = 16'b0000010111000000;
            15'd28077: log10_cal = 16'b0000010111000000;
            15'd28078: log10_cal = 16'b0000010111000000;
            15'd28079: log10_cal = 16'b0000010111000000;
            15'd28080: log10_cal = 16'b0000010111000000;
            15'd28081: log10_cal = 16'b0000010111000000;
            15'd28082: log10_cal = 16'b0000010111000000;
            15'd28083: log10_cal = 16'b0000010111000000;
            15'd28084: log10_cal = 16'b0000010111000000;
            15'd28085: log10_cal = 16'b0000010111000000;
            15'd28086: log10_cal = 16'b0000010111000000;
            15'd28087: log10_cal = 16'b0000010111000000;
            15'd28088: log10_cal = 16'b0000010111000000;
            15'd28089: log10_cal = 16'b0000010111000000;
            15'd28090: log10_cal = 16'b0000010111000000;
            15'd28091: log10_cal = 16'b0000010111000000;
            15'd28092: log10_cal = 16'b0000010111000000;
            15'd28093: log10_cal = 16'b0000010111000000;
            15'd28094: log10_cal = 16'b0000010111000000;
            15'd28095: log10_cal = 16'b0000010111000000;
            15'd28096: log10_cal = 16'b0000010111000000;
            15'd28097: log10_cal = 16'b0000010111000000;
            15'd28098: log10_cal = 16'b0000010111000000;
            15'd28099: log10_cal = 16'b0000010111000000;
            15'd28100: log10_cal = 16'b0000010111000000;
            15'd28101: log10_cal = 16'b0000010111000000;
            15'd28102: log10_cal = 16'b0000010111000000;
            15'd28103: log10_cal = 16'b0000010111000000;
            15'd28104: log10_cal = 16'b0000010111000000;
            15'd28105: log10_cal = 16'b0000010111000001;
            15'd28106: log10_cal = 16'b0000010111000001;
            15'd28107: log10_cal = 16'b0000010111000001;
            15'd28108: log10_cal = 16'b0000010111000001;
            15'd28109: log10_cal = 16'b0000010111000001;
            15'd28110: log10_cal = 16'b0000010111000001;
            15'd28111: log10_cal = 16'b0000010111000001;
            15'd28112: log10_cal = 16'b0000010111000001;
            15'd28113: log10_cal = 16'b0000010111000001;
            15'd28114: log10_cal = 16'b0000010111000001;
            15'd28115: log10_cal = 16'b0000010111000001;
            15'd28116: log10_cal = 16'b0000010111000001;
            15'd28117: log10_cal = 16'b0000010111000001;
            15'd28118: log10_cal = 16'b0000010111000001;
            15'd28119: log10_cal = 16'b0000010111000001;
            15'd28120: log10_cal = 16'b0000010111000001;
            15'd28121: log10_cal = 16'b0000010111000001;
            15'd28122: log10_cal = 16'b0000010111000001;
            15'd28123: log10_cal = 16'b0000010111000001;
            15'd28124: log10_cal = 16'b0000010111000001;
            15'd28125: log10_cal = 16'b0000010111000001;
            15'd28126: log10_cal = 16'b0000010111000001;
            15'd28127: log10_cal = 16'b0000010111000001;
            15'd28128: log10_cal = 16'b0000010111000001;
            15'd28129: log10_cal = 16'b0000010111000001;
            15'd28130: log10_cal = 16'b0000010111000001;
            15'd28131: log10_cal = 16'b0000010111000001;
            15'd28132: log10_cal = 16'b0000010111000001;
            15'd28133: log10_cal = 16'b0000010111000001;
            15'd28134: log10_cal = 16'b0000010111000001;
            15'd28135: log10_cal = 16'b0000010111000001;
            15'd28136: log10_cal = 16'b0000010111000001;
            15'd28137: log10_cal = 16'b0000010111000001;
            15'd28138: log10_cal = 16'b0000010111000001;
            15'd28139: log10_cal = 16'b0000010111000001;
            15'd28140: log10_cal = 16'b0000010111000001;
            15'd28141: log10_cal = 16'b0000010111000001;
            15'd28142: log10_cal = 16'b0000010111000001;
            15'd28143: log10_cal = 16'b0000010111000001;
            15'd28144: log10_cal = 16'b0000010111000001;
            15'd28145: log10_cal = 16'b0000010111000001;
            15'd28146: log10_cal = 16'b0000010111000001;
            15'd28147: log10_cal = 16'b0000010111000001;
            15'd28148: log10_cal = 16'b0000010111000001;
            15'd28149: log10_cal = 16'b0000010111000001;
            15'd28150: log10_cal = 16'b0000010111000001;
            15'd28151: log10_cal = 16'b0000010111000001;
            15'd28152: log10_cal = 16'b0000010111000001;
            15'd28153: log10_cal = 16'b0000010111000001;
            15'd28154: log10_cal = 16'b0000010111000001;
            15'd28155: log10_cal = 16'b0000010111000001;
            15'd28156: log10_cal = 16'b0000010111000001;
            15'd28157: log10_cal = 16'b0000010111000001;
            15'd28158: log10_cal = 16'b0000010111000001;
            15'd28159: log10_cal = 16'b0000010111000001;
            15'd28160: log10_cal = 16'b0000010111000001;
            15'd28161: log10_cal = 16'b0000010111000001;
            15'd28162: log10_cal = 16'b0000010111000001;
            15'd28163: log10_cal = 16'b0000010111000001;
            15'd28164: log10_cal = 16'b0000010111000001;
            15'd28165: log10_cal = 16'b0000010111000001;
            15'd28166: log10_cal = 16'b0000010111000001;
            15'd28167: log10_cal = 16'b0000010111000001;
            15'd28168: log10_cal = 16'b0000010111000010;
            15'd28169: log10_cal = 16'b0000010111000010;
            15'd28170: log10_cal = 16'b0000010111000010;
            15'd28171: log10_cal = 16'b0000010111000010;
            15'd28172: log10_cal = 16'b0000010111000010;
            15'd28173: log10_cal = 16'b0000010111000010;
            15'd28174: log10_cal = 16'b0000010111000010;
            15'd28175: log10_cal = 16'b0000010111000010;
            15'd28176: log10_cal = 16'b0000010111000010;
            15'd28177: log10_cal = 16'b0000010111000010;
            15'd28178: log10_cal = 16'b0000010111000010;
            15'd28179: log10_cal = 16'b0000010111000010;
            15'd28180: log10_cal = 16'b0000010111000010;
            15'd28181: log10_cal = 16'b0000010111000010;
            15'd28182: log10_cal = 16'b0000010111000010;
            15'd28183: log10_cal = 16'b0000010111000010;
            15'd28184: log10_cal = 16'b0000010111000010;
            15'd28185: log10_cal = 16'b0000010111000010;
            15'd28186: log10_cal = 16'b0000010111000010;
            15'd28187: log10_cal = 16'b0000010111000010;
            15'd28188: log10_cal = 16'b0000010111000010;
            15'd28189: log10_cal = 16'b0000010111000010;
            15'd28190: log10_cal = 16'b0000010111000010;
            15'd28191: log10_cal = 16'b0000010111000010;
            15'd28192: log10_cal = 16'b0000010111000010;
            15'd28193: log10_cal = 16'b0000010111000010;
            15'd28194: log10_cal = 16'b0000010111000010;
            15'd28195: log10_cal = 16'b0000010111000010;
            15'd28196: log10_cal = 16'b0000010111000010;
            15'd28197: log10_cal = 16'b0000010111000010;
            15'd28198: log10_cal = 16'b0000010111000010;
            15'd28199: log10_cal = 16'b0000010111000010;
            15'd28200: log10_cal = 16'b0000010111000010;
            15'd28201: log10_cal = 16'b0000010111000010;
            15'd28202: log10_cal = 16'b0000010111000010;
            15'd28203: log10_cal = 16'b0000010111000010;
            15'd28204: log10_cal = 16'b0000010111000010;
            15'd28205: log10_cal = 16'b0000010111000010;
            15'd28206: log10_cal = 16'b0000010111000010;
            15'd28207: log10_cal = 16'b0000010111000010;
            15'd28208: log10_cal = 16'b0000010111000010;
            15'd28209: log10_cal = 16'b0000010111000010;
            15'd28210: log10_cal = 16'b0000010111000010;
            15'd28211: log10_cal = 16'b0000010111000010;
            15'd28212: log10_cal = 16'b0000010111000010;
            15'd28213: log10_cal = 16'b0000010111000010;
            15'd28214: log10_cal = 16'b0000010111000010;
            15'd28215: log10_cal = 16'b0000010111000010;
            15'd28216: log10_cal = 16'b0000010111000010;
            15'd28217: log10_cal = 16'b0000010111000010;
            15'd28218: log10_cal = 16'b0000010111000010;
            15'd28219: log10_cal = 16'b0000010111000010;
            15'd28220: log10_cal = 16'b0000010111000010;
            15'd28221: log10_cal = 16'b0000010111000010;
            15'd28222: log10_cal = 16'b0000010111000010;
            15'd28223: log10_cal = 16'b0000010111000010;
            15'd28224: log10_cal = 16'b0000010111000010;
            15'd28225: log10_cal = 16'b0000010111000010;
            15'd28226: log10_cal = 16'b0000010111000010;
            15'd28227: log10_cal = 16'b0000010111000010;
            15'd28228: log10_cal = 16'b0000010111000010;
            15'd28229: log10_cal = 16'b0000010111000010;
            15'd28230: log10_cal = 16'b0000010111000010;
            15'd28231: log10_cal = 16'b0000010111000010;
            15'd28232: log10_cal = 16'b0000010111000011;
            15'd28233: log10_cal = 16'b0000010111000011;
            15'd28234: log10_cal = 16'b0000010111000011;
            15'd28235: log10_cal = 16'b0000010111000011;
            15'd28236: log10_cal = 16'b0000010111000011;
            15'd28237: log10_cal = 16'b0000010111000011;
            15'd28238: log10_cal = 16'b0000010111000011;
            15'd28239: log10_cal = 16'b0000010111000011;
            15'd28240: log10_cal = 16'b0000010111000011;
            15'd28241: log10_cal = 16'b0000010111000011;
            15'd28242: log10_cal = 16'b0000010111000011;
            15'd28243: log10_cal = 16'b0000010111000011;
            15'd28244: log10_cal = 16'b0000010111000011;
            15'd28245: log10_cal = 16'b0000010111000011;
            15'd28246: log10_cal = 16'b0000010111000011;
            15'd28247: log10_cal = 16'b0000010111000011;
            15'd28248: log10_cal = 16'b0000010111000011;
            15'd28249: log10_cal = 16'b0000010111000011;
            15'd28250: log10_cal = 16'b0000010111000011;
            15'd28251: log10_cal = 16'b0000010111000011;
            15'd28252: log10_cal = 16'b0000010111000011;
            15'd28253: log10_cal = 16'b0000010111000011;
            15'd28254: log10_cal = 16'b0000010111000011;
            15'd28255: log10_cal = 16'b0000010111000011;
            15'd28256: log10_cal = 16'b0000010111000011;
            15'd28257: log10_cal = 16'b0000010111000011;
            15'd28258: log10_cal = 16'b0000010111000011;
            15'd28259: log10_cal = 16'b0000010111000011;
            15'd28260: log10_cal = 16'b0000010111000011;
            15'd28261: log10_cal = 16'b0000010111000011;
            15'd28262: log10_cal = 16'b0000010111000011;
            15'd28263: log10_cal = 16'b0000010111000011;
            15'd28264: log10_cal = 16'b0000010111000011;
            15'd28265: log10_cal = 16'b0000010111000011;
            15'd28266: log10_cal = 16'b0000010111000011;
            15'd28267: log10_cal = 16'b0000010111000011;
            15'd28268: log10_cal = 16'b0000010111000011;
            15'd28269: log10_cal = 16'b0000010111000011;
            15'd28270: log10_cal = 16'b0000010111000011;
            15'd28271: log10_cal = 16'b0000010111000011;
            15'd28272: log10_cal = 16'b0000010111000011;
            15'd28273: log10_cal = 16'b0000010111000011;
            15'd28274: log10_cal = 16'b0000010111000011;
            15'd28275: log10_cal = 16'b0000010111000011;
            15'd28276: log10_cal = 16'b0000010111000011;
            15'd28277: log10_cal = 16'b0000010111000011;
            15'd28278: log10_cal = 16'b0000010111000011;
            15'd28279: log10_cal = 16'b0000010111000011;
            15'd28280: log10_cal = 16'b0000010111000011;
            15'd28281: log10_cal = 16'b0000010111000011;
            15'd28282: log10_cal = 16'b0000010111000011;
            15'd28283: log10_cal = 16'b0000010111000011;
            15'd28284: log10_cal = 16'b0000010111000011;
            15'd28285: log10_cal = 16'b0000010111000011;
            15'd28286: log10_cal = 16'b0000010111000011;
            15'd28287: log10_cal = 16'b0000010111000011;
            15'd28288: log10_cal = 16'b0000010111000011;
            15'd28289: log10_cal = 16'b0000010111000011;
            15'd28290: log10_cal = 16'b0000010111000011;
            15'd28291: log10_cal = 16'b0000010111000011;
            15'd28292: log10_cal = 16'b0000010111000011;
            15'd28293: log10_cal = 16'b0000010111000011;
            15'd28294: log10_cal = 16'b0000010111000011;
            15'd28295: log10_cal = 16'b0000010111000100;
            15'd28296: log10_cal = 16'b0000010111000100;
            15'd28297: log10_cal = 16'b0000010111000100;
            15'd28298: log10_cal = 16'b0000010111000100;
            15'd28299: log10_cal = 16'b0000010111000100;
            15'd28300: log10_cal = 16'b0000010111000100;
            15'd28301: log10_cal = 16'b0000010111000100;
            15'd28302: log10_cal = 16'b0000010111000100;
            15'd28303: log10_cal = 16'b0000010111000100;
            15'd28304: log10_cal = 16'b0000010111000100;
            15'd28305: log10_cal = 16'b0000010111000100;
            15'd28306: log10_cal = 16'b0000010111000100;
            15'd28307: log10_cal = 16'b0000010111000100;
            15'd28308: log10_cal = 16'b0000010111000100;
            15'd28309: log10_cal = 16'b0000010111000100;
            15'd28310: log10_cal = 16'b0000010111000100;
            15'd28311: log10_cal = 16'b0000010111000100;
            15'd28312: log10_cal = 16'b0000010111000100;
            15'd28313: log10_cal = 16'b0000010111000100;
            15'd28314: log10_cal = 16'b0000010111000100;
            15'd28315: log10_cal = 16'b0000010111000100;
            15'd28316: log10_cal = 16'b0000010111000100;
            15'd28317: log10_cal = 16'b0000010111000100;
            15'd28318: log10_cal = 16'b0000010111000100;
            15'd28319: log10_cal = 16'b0000010111000100;
            15'd28320: log10_cal = 16'b0000010111000100;
            15'd28321: log10_cal = 16'b0000010111000100;
            15'd28322: log10_cal = 16'b0000010111000100;
            15'd28323: log10_cal = 16'b0000010111000100;
            15'd28324: log10_cal = 16'b0000010111000100;
            15'd28325: log10_cal = 16'b0000010111000100;
            15'd28326: log10_cal = 16'b0000010111000100;
            15'd28327: log10_cal = 16'b0000010111000100;
            15'd28328: log10_cal = 16'b0000010111000100;
            15'd28329: log10_cal = 16'b0000010111000100;
            15'd28330: log10_cal = 16'b0000010111000100;
            15'd28331: log10_cal = 16'b0000010111000100;
            15'd28332: log10_cal = 16'b0000010111000100;
            15'd28333: log10_cal = 16'b0000010111000100;
            15'd28334: log10_cal = 16'b0000010111000100;
            15'd28335: log10_cal = 16'b0000010111000100;
            15'd28336: log10_cal = 16'b0000010111000100;
            15'd28337: log10_cal = 16'b0000010111000100;
            15'd28338: log10_cal = 16'b0000010111000100;
            15'd28339: log10_cal = 16'b0000010111000100;
            15'd28340: log10_cal = 16'b0000010111000100;
            15'd28341: log10_cal = 16'b0000010111000100;
            15'd28342: log10_cal = 16'b0000010111000100;
            15'd28343: log10_cal = 16'b0000010111000100;
            15'd28344: log10_cal = 16'b0000010111000100;
            15'd28345: log10_cal = 16'b0000010111000100;
            15'd28346: log10_cal = 16'b0000010111000100;
            15'd28347: log10_cal = 16'b0000010111000100;
            15'd28348: log10_cal = 16'b0000010111000100;
            15'd28349: log10_cal = 16'b0000010111000100;
            15'd28350: log10_cal = 16'b0000010111000100;
            15'd28351: log10_cal = 16'b0000010111000100;
            15'd28352: log10_cal = 16'b0000010111000100;
            15'd28353: log10_cal = 16'b0000010111000100;
            15'd28354: log10_cal = 16'b0000010111000100;
            15'd28355: log10_cal = 16'b0000010111000100;
            15'd28356: log10_cal = 16'b0000010111000100;
            15'd28357: log10_cal = 16'b0000010111000100;
            15'd28358: log10_cal = 16'b0000010111000100;
            15'd28359: log10_cal = 16'b0000010111000101;
            15'd28360: log10_cal = 16'b0000010111000101;
            15'd28361: log10_cal = 16'b0000010111000101;
            15'd28362: log10_cal = 16'b0000010111000101;
            15'd28363: log10_cal = 16'b0000010111000101;
            15'd28364: log10_cal = 16'b0000010111000101;
            15'd28365: log10_cal = 16'b0000010111000101;
            15'd28366: log10_cal = 16'b0000010111000101;
            15'd28367: log10_cal = 16'b0000010111000101;
            15'd28368: log10_cal = 16'b0000010111000101;
            15'd28369: log10_cal = 16'b0000010111000101;
            15'd28370: log10_cal = 16'b0000010111000101;
            15'd28371: log10_cal = 16'b0000010111000101;
            15'd28372: log10_cal = 16'b0000010111000101;
            15'd28373: log10_cal = 16'b0000010111000101;
            15'd28374: log10_cal = 16'b0000010111000101;
            15'd28375: log10_cal = 16'b0000010111000101;
            15'd28376: log10_cal = 16'b0000010111000101;
            15'd28377: log10_cal = 16'b0000010111000101;
            15'd28378: log10_cal = 16'b0000010111000101;
            15'd28379: log10_cal = 16'b0000010111000101;
            15'd28380: log10_cal = 16'b0000010111000101;
            15'd28381: log10_cal = 16'b0000010111000101;
            15'd28382: log10_cal = 16'b0000010111000101;
            15'd28383: log10_cal = 16'b0000010111000101;
            15'd28384: log10_cal = 16'b0000010111000101;
            15'd28385: log10_cal = 16'b0000010111000101;
            15'd28386: log10_cal = 16'b0000010111000101;
            15'd28387: log10_cal = 16'b0000010111000101;
            15'd28388: log10_cal = 16'b0000010111000101;
            15'd28389: log10_cal = 16'b0000010111000101;
            15'd28390: log10_cal = 16'b0000010111000101;
            15'd28391: log10_cal = 16'b0000010111000101;
            15'd28392: log10_cal = 16'b0000010111000101;
            15'd28393: log10_cal = 16'b0000010111000101;
            15'd28394: log10_cal = 16'b0000010111000101;
            15'd28395: log10_cal = 16'b0000010111000101;
            15'd28396: log10_cal = 16'b0000010111000101;
            15'd28397: log10_cal = 16'b0000010111000101;
            15'd28398: log10_cal = 16'b0000010111000101;
            15'd28399: log10_cal = 16'b0000010111000101;
            15'd28400: log10_cal = 16'b0000010111000101;
            15'd28401: log10_cal = 16'b0000010111000101;
            15'd28402: log10_cal = 16'b0000010111000101;
            15'd28403: log10_cal = 16'b0000010111000101;
            15'd28404: log10_cal = 16'b0000010111000101;
            15'd28405: log10_cal = 16'b0000010111000101;
            15'd28406: log10_cal = 16'b0000010111000101;
            15'd28407: log10_cal = 16'b0000010111000101;
            15'd28408: log10_cal = 16'b0000010111000101;
            15'd28409: log10_cal = 16'b0000010111000101;
            15'd28410: log10_cal = 16'b0000010111000101;
            15'd28411: log10_cal = 16'b0000010111000101;
            15'd28412: log10_cal = 16'b0000010111000101;
            15'd28413: log10_cal = 16'b0000010111000101;
            15'd28414: log10_cal = 16'b0000010111000101;
            15'd28415: log10_cal = 16'b0000010111000101;
            15'd28416: log10_cal = 16'b0000010111000101;
            15'd28417: log10_cal = 16'b0000010111000101;
            15'd28418: log10_cal = 16'b0000010111000101;
            15'd28419: log10_cal = 16'b0000010111000101;
            15'd28420: log10_cal = 16'b0000010111000101;
            15'd28421: log10_cal = 16'b0000010111000101;
            15'd28422: log10_cal = 16'b0000010111000101;
            15'd28423: log10_cal = 16'b0000010111000110;
            15'd28424: log10_cal = 16'b0000010111000110;
            15'd28425: log10_cal = 16'b0000010111000110;
            15'd28426: log10_cal = 16'b0000010111000110;
            15'd28427: log10_cal = 16'b0000010111000110;
            15'd28428: log10_cal = 16'b0000010111000110;
            15'd28429: log10_cal = 16'b0000010111000110;
            15'd28430: log10_cal = 16'b0000010111000110;
            15'd28431: log10_cal = 16'b0000010111000110;
            15'd28432: log10_cal = 16'b0000010111000110;
            15'd28433: log10_cal = 16'b0000010111000110;
            15'd28434: log10_cal = 16'b0000010111000110;
            15'd28435: log10_cal = 16'b0000010111000110;
            15'd28436: log10_cal = 16'b0000010111000110;
            15'd28437: log10_cal = 16'b0000010111000110;
            15'd28438: log10_cal = 16'b0000010111000110;
            15'd28439: log10_cal = 16'b0000010111000110;
            15'd28440: log10_cal = 16'b0000010111000110;
            15'd28441: log10_cal = 16'b0000010111000110;
            15'd28442: log10_cal = 16'b0000010111000110;
            15'd28443: log10_cal = 16'b0000010111000110;
            15'd28444: log10_cal = 16'b0000010111000110;
            15'd28445: log10_cal = 16'b0000010111000110;
            15'd28446: log10_cal = 16'b0000010111000110;
            15'd28447: log10_cal = 16'b0000010111000110;
            15'd28448: log10_cal = 16'b0000010111000110;
            15'd28449: log10_cal = 16'b0000010111000110;
            15'd28450: log10_cal = 16'b0000010111000110;
            15'd28451: log10_cal = 16'b0000010111000110;
            15'd28452: log10_cal = 16'b0000010111000110;
            15'd28453: log10_cal = 16'b0000010111000110;
            15'd28454: log10_cal = 16'b0000010111000110;
            15'd28455: log10_cal = 16'b0000010111000110;
            15'd28456: log10_cal = 16'b0000010111000110;
            15'd28457: log10_cal = 16'b0000010111000110;
            15'd28458: log10_cal = 16'b0000010111000110;
            15'd28459: log10_cal = 16'b0000010111000110;
            15'd28460: log10_cal = 16'b0000010111000110;
            15'd28461: log10_cal = 16'b0000010111000110;
            15'd28462: log10_cal = 16'b0000010111000110;
            15'd28463: log10_cal = 16'b0000010111000110;
            15'd28464: log10_cal = 16'b0000010111000110;
            15'd28465: log10_cal = 16'b0000010111000110;
            15'd28466: log10_cal = 16'b0000010111000110;
            15'd28467: log10_cal = 16'b0000010111000110;
            15'd28468: log10_cal = 16'b0000010111000110;
            15'd28469: log10_cal = 16'b0000010111000110;
            15'd28470: log10_cal = 16'b0000010111000110;
            15'd28471: log10_cal = 16'b0000010111000110;
            15'd28472: log10_cal = 16'b0000010111000110;
            15'd28473: log10_cal = 16'b0000010111000110;
            15'd28474: log10_cal = 16'b0000010111000110;
            15'd28475: log10_cal = 16'b0000010111000110;
            15'd28476: log10_cal = 16'b0000010111000110;
            15'd28477: log10_cal = 16'b0000010111000110;
            15'd28478: log10_cal = 16'b0000010111000110;
            15'd28479: log10_cal = 16'b0000010111000110;
            15'd28480: log10_cal = 16'b0000010111000110;
            15'd28481: log10_cal = 16'b0000010111000110;
            15'd28482: log10_cal = 16'b0000010111000110;
            15'd28483: log10_cal = 16'b0000010111000110;
            15'd28484: log10_cal = 16'b0000010111000110;
            15'd28485: log10_cal = 16'b0000010111000110;
            15'd28486: log10_cal = 16'b0000010111000110;
            15'd28487: log10_cal = 16'b0000010111000111;
            15'd28488: log10_cal = 16'b0000010111000111;
            15'd28489: log10_cal = 16'b0000010111000111;
            15'd28490: log10_cal = 16'b0000010111000111;
            15'd28491: log10_cal = 16'b0000010111000111;
            15'd28492: log10_cal = 16'b0000010111000111;
            15'd28493: log10_cal = 16'b0000010111000111;
            15'd28494: log10_cal = 16'b0000010111000111;
            15'd28495: log10_cal = 16'b0000010111000111;
            15'd28496: log10_cal = 16'b0000010111000111;
            15'd28497: log10_cal = 16'b0000010111000111;
            15'd28498: log10_cal = 16'b0000010111000111;
            15'd28499: log10_cal = 16'b0000010111000111;
            15'd28500: log10_cal = 16'b0000010111000111;
            15'd28501: log10_cal = 16'b0000010111000111;
            15'd28502: log10_cal = 16'b0000010111000111;
            15'd28503: log10_cal = 16'b0000010111000111;
            15'd28504: log10_cal = 16'b0000010111000111;
            15'd28505: log10_cal = 16'b0000010111000111;
            15'd28506: log10_cal = 16'b0000010111000111;
            15'd28507: log10_cal = 16'b0000010111000111;
            15'd28508: log10_cal = 16'b0000010111000111;
            15'd28509: log10_cal = 16'b0000010111000111;
            15'd28510: log10_cal = 16'b0000010111000111;
            15'd28511: log10_cal = 16'b0000010111000111;
            15'd28512: log10_cal = 16'b0000010111000111;
            15'd28513: log10_cal = 16'b0000010111000111;
            15'd28514: log10_cal = 16'b0000010111000111;
            15'd28515: log10_cal = 16'b0000010111000111;
            15'd28516: log10_cal = 16'b0000010111000111;
            15'd28517: log10_cal = 16'b0000010111000111;
            15'd28518: log10_cal = 16'b0000010111000111;
            15'd28519: log10_cal = 16'b0000010111000111;
            15'd28520: log10_cal = 16'b0000010111000111;
            15'd28521: log10_cal = 16'b0000010111000111;
            15'd28522: log10_cal = 16'b0000010111000111;
            15'd28523: log10_cal = 16'b0000010111000111;
            15'd28524: log10_cal = 16'b0000010111000111;
            15'd28525: log10_cal = 16'b0000010111000111;
            15'd28526: log10_cal = 16'b0000010111000111;
            15'd28527: log10_cal = 16'b0000010111000111;
            15'd28528: log10_cal = 16'b0000010111000111;
            15'd28529: log10_cal = 16'b0000010111000111;
            15'd28530: log10_cal = 16'b0000010111000111;
            15'd28531: log10_cal = 16'b0000010111000111;
            15'd28532: log10_cal = 16'b0000010111000111;
            15'd28533: log10_cal = 16'b0000010111000111;
            15'd28534: log10_cal = 16'b0000010111000111;
            15'd28535: log10_cal = 16'b0000010111000111;
            15'd28536: log10_cal = 16'b0000010111000111;
            15'd28537: log10_cal = 16'b0000010111000111;
            15'd28538: log10_cal = 16'b0000010111000111;
            15'd28539: log10_cal = 16'b0000010111000111;
            15'd28540: log10_cal = 16'b0000010111000111;
            15'd28541: log10_cal = 16'b0000010111000111;
            15'd28542: log10_cal = 16'b0000010111000111;
            15'd28543: log10_cal = 16'b0000010111000111;
            15'd28544: log10_cal = 16'b0000010111000111;
            15'd28545: log10_cal = 16'b0000010111000111;
            15'd28546: log10_cal = 16'b0000010111000111;
            15'd28547: log10_cal = 16'b0000010111000111;
            15'd28548: log10_cal = 16'b0000010111000111;
            15'd28549: log10_cal = 16'b0000010111000111;
            15'd28550: log10_cal = 16'b0000010111000111;
            15'd28551: log10_cal = 16'b0000010111001000;
            15'd28552: log10_cal = 16'b0000010111001000;
            15'd28553: log10_cal = 16'b0000010111001000;
            15'd28554: log10_cal = 16'b0000010111001000;
            15'd28555: log10_cal = 16'b0000010111001000;
            15'd28556: log10_cal = 16'b0000010111001000;
            15'd28557: log10_cal = 16'b0000010111001000;
            15'd28558: log10_cal = 16'b0000010111001000;
            15'd28559: log10_cal = 16'b0000010111001000;
            15'd28560: log10_cal = 16'b0000010111001000;
            15'd28561: log10_cal = 16'b0000010111001000;
            15'd28562: log10_cal = 16'b0000010111001000;
            15'd28563: log10_cal = 16'b0000010111001000;
            15'd28564: log10_cal = 16'b0000010111001000;
            15'd28565: log10_cal = 16'b0000010111001000;
            15'd28566: log10_cal = 16'b0000010111001000;
            15'd28567: log10_cal = 16'b0000010111001000;
            15'd28568: log10_cal = 16'b0000010111001000;
            15'd28569: log10_cal = 16'b0000010111001000;
            15'd28570: log10_cal = 16'b0000010111001000;
            15'd28571: log10_cal = 16'b0000010111001000;
            15'd28572: log10_cal = 16'b0000010111001000;
            15'd28573: log10_cal = 16'b0000010111001000;
            15'd28574: log10_cal = 16'b0000010111001000;
            15'd28575: log10_cal = 16'b0000010111001000;
            15'd28576: log10_cal = 16'b0000010111001000;
            15'd28577: log10_cal = 16'b0000010111001000;
            15'd28578: log10_cal = 16'b0000010111001000;
            15'd28579: log10_cal = 16'b0000010111001000;
            15'd28580: log10_cal = 16'b0000010111001000;
            15'd28581: log10_cal = 16'b0000010111001000;
            15'd28582: log10_cal = 16'b0000010111001000;
            15'd28583: log10_cal = 16'b0000010111001000;
            15'd28584: log10_cal = 16'b0000010111001000;
            15'd28585: log10_cal = 16'b0000010111001000;
            15'd28586: log10_cal = 16'b0000010111001000;
            15'd28587: log10_cal = 16'b0000010111001000;
            15'd28588: log10_cal = 16'b0000010111001000;
            15'd28589: log10_cal = 16'b0000010111001000;
            15'd28590: log10_cal = 16'b0000010111001000;
            15'd28591: log10_cal = 16'b0000010111001000;
            15'd28592: log10_cal = 16'b0000010111001000;
            15'd28593: log10_cal = 16'b0000010111001000;
            15'd28594: log10_cal = 16'b0000010111001000;
            15'd28595: log10_cal = 16'b0000010111001000;
            15'd28596: log10_cal = 16'b0000010111001000;
            15'd28597: log10_cal = 16'b0000010111001000;
            15'd28598: log10_cal = 16'b0000010111001000;
            15'd28599: log10_cal = 16'b0000010111001000;
            15'd28600: log10_cal = 16'b0000010111001000;
            15'd28601: log10_cal = 16'b0000010111001000;
            15'd28602: log10_cal = 16'b0000010111001000;
            15'd28603: log10_cal = 16'b0000010111001000;
            15'd28604: log10_cal = 16'b0000010111001000;
            15'd28605: log10_cal = 16'b0000010111001000;
            15'd28606: log10_cal = 16'b0000010111001000;
            15'd28607: log10_cal = 16'b0000010111001000;
            15'd28608: log10_cal = 16'b0000010111001000;
            15'd28609: log10_cal = 16'b0000010111001000;
            15'd28610: log10_cal = 16'b0000010111001000;
            15'd28611: log10_cal = 16'b0000010111001000;
            15'd28612: log10_cal = 16'b0000010111001000;
            15'd28613: log10_cal = 16'b0000010111001000;
            15'd28614: log10_cal = 16'b0000010111001000;
            15'd28615: log10_cal = 16'b0000010111001001;
            15'd28616: log10_cal = 16'b0000010111001001;
            15'd28617: log10_cal = 16'b0000010111001001;
            15'd28618: log10_cal = 16'b0000010111001001;
            15'd28619: log10_cal = 16'b0000010111001001;
            15'd28620: log10_cal = 16'b0000010111001001;
            15'd28621: log10_cal = 16'b0000010111001001;
            15'd28622: log10_cal = 16'b0000010111001001;
            15'd28623: log10_cal = 16'b0000010111001001;
            15'd28624: log10_cal = 16'b0000010111001001;
            15'd28625: log10_cal = 16'b0000010111001001;
            15'd28626: log10_cal = 16'b0000010111001001;
            15'd28627: log10_cal = 16'b0000010111001001;
            15'd28628: log10_cal = 16'b0000010111001001;
            15'd28629: log10_cal = 16'b0000010111001001;
            15'd28630: log10_cal = 16'b0000010111001001;
            15'd28631: log10_cal = 16'b0000010111001001;
            15'd28632: log10_cal = 16'b0000010111001001;
            15'd28633: log10_cal = 16'b0000010111001001;
            15'd28634: log10_cal = 16'b0000010111001001;
            15'd28635: log10_cal = 16'b0000010111001001;
            15'd28636: log10_cal = 16'b0000010111001001;
            15'd28637: log10_cal = 16'b0000010111001001;
            15'd28638: log10_cal = 16'b0000010111001001;
            15'd28639: log10_cal = 16'b0000010111001001;
            15'd28640: log10_cal = 16'b0000010111001001;
            15'd28641: log10_cal = 16'b0000010111001001;
            15'd28642: log10_cal = 16'b0000010111001001;
            15'd28643: log10_cal = 16'b0000010111001001;
            15'd28644: log10_cal = 16'b0000010111001001;
            15'd28645: log10_cal = 16'b0000010111001001;
            15'd28646: log10_cal = 16'b0000010111001001;
            15'd28647: log10_cal = 16'b0000010111001001;
            15'd28648: log10_cal = 16'b0000010111001001;
            15'd28649: log10_cal = 16'b0000010111001001;
            15'd28650: log10_cal = 16'b0000010111001001;
            15'd28651: log10_cal = 16'b0000010111001001;
            15'd28652: log10_cal = 16'b0000010111001001;
            15'd28653: log10_cal = 16'b0000010111001001;
            15'd28654: log10_cal = 16'b0000010111001001;
            15'd28655: log10_cal = 16'b0000010111001001;
            15'd28656: log10_cal = 16'b0000010111001001;
            15'd28657: log10_cal = 16'b0000010111001001;
            15'd28658: log10_cal = 16'b0000010111001001;
            15'd28659: log10_cal = 16'b0000010111001001;
            15'd28660: log10_cal = 16'b0000010111001001;
            15'd28661: log10_cal = 16'b0000010111001001;
            15'd28662: log10_cal = 16'b0000010111001001;
            15'd28663: log10_cal = 16'b0000010111001001;
            15'd28664: log10_cal = 16'b0000010111001001;
            15'd28665: log10_cal = 16'b0000010111001001;
            15'd28666: log10_cal = 16'b0000010111001001;
            15'd28667: log10_cal = 16'b0000010111001001;
            15'd28668: log10_cal = 16'b0000010111001001;
            15'd28669: log10_cal = 16'b0000010111001001;
            15'd28670: log10_cal = 16'b0000010111001001;
            15'd28671: log10_cal = 16'b0000010111001001;
            15'd28672: log10_cal = 16'b0000010111001001;
            15'd28673: log10_cal = 16'b0000010111001001;
            15'd28674: log10_cal = 16'b0000010111001001;
            15'd28675: log10_cal = 16'b0000010111001001;
            15'd28676: log10_cal = 16'b0000010111001001;
            15'd28677: log10_cal = 16'b0000010111001001;
            15'd28678: log10_cal = 16'b0000010111001001;
            15'd28679: log10_cal = 16'b0000010111001001;
            15'd28680: log10_cal = 16'b0000010111001010;
            15'd28681: log10_cal = 16'b0000010111001010;
            15'd28682: log10_cal = 16'b0000010111001010;
            15'd28683: log10_cal = 16'b0000010111001010;
            15'd28684: log10_cal = 16'b0000010111001010;
            15'd28685: log10_cal = 16'b0000010111001010;
            15'd28686: log10_cal = 16'b0000010111001010;
            15'd28687: log10_cal = 16'b0000010111001010;
            15'd28688: log10_cal = 16'b0000010111001010;
            15'd28689: log10_cal = 16'b0000010111001010;
            15'd28690: log10_cal = 16'b0000010111001010;
            15'd28691: log10_cal = 16'b0000010111001010;
            15'd28692: log10_cal = 16'b0000010111001010;
            15'd28693: log10_cal = 16'b0000010111001010;
            15'd28694: log10_cal = 16'b0000010111001010;
            15'd28695: log10_cal = 16'b0000010111001010;
            15'd28696: log10_cal = 16'b0000010111001010;
            15'd28697: log10_cal = 16'b0000010111001010;
            15'd28698: log10_cal = 16'b0000010111001010;
            15'd28699: log10_cal = 16'b0000010111001010;
            15'd28700: log10_cal = 16'b0000010111001010;
            15'd28701: log10_cal = 16'b0000010111001010;
            15'd28702: log10_cal = 16'b0000010111001010;
            15'd28703: log10_cal = 16'b0000010111001010;
            15'd28704: log10_cal = 16'b0000010111001010;
            15'd28705: log10_cal = 16'b0000010111001010;
            15'd28706: log10_cal = 16'b0000010111001010;
            15'd28707: log10_cal = 16'b0000010111001010;
            15'd28708: log10_cal = 16'b0000010111001010;
            15'd28709: log10_cal = 16'b0000010111001010;
            15'd28710: log10_cal = 16'b0000010111001010;
            15'd28711: log10_cal = 16'b0000010111001010;
            15'd28712: log10_cal = 16'b0000010111001010;
            15'd28713: log10_cal = 16'b0000010111001010;
            15'd28714: log10_cal = 16'b0000010111001010;
            15'd28715: log10_cal = 16'b0000010111001010;
            15'd28716: log10_cal = 16'b0000010111001010;
            15'd28717: log10_cal = 16'b0000010111001010;
            15'd28718: log10_cal = 16'b0000010111001010;
            15'd28719: log10_cal = 16'b0000010111001010;
            15'd28720: log10_cal = 16'b0000010111001010;
            15'd28721: log10_cal = 16'b0000010111001010;
            15'd28722: log10_cal = 16'b0000010111001010;
            15'd28723: log10_cal = 16'b0000010111001010;
            15'd28724: log10_cal = 16'b0000010111001010;
            15'd28725: log10_cal = 16'b0000010111001010;
            15'd28726: log10_cal = 16'b0000010111001010;
            15'd28727: log10_cal = 16'b0000010111001010;
            15'd28728: log10_cal = 16'b0000010111001010;
            15'd28729: log10_cal = 16'b0000010111001010;
            15'd28730: log10_cal = 16'b0000010111001010;
            15'd28731: log10_cal = 16'b0000010111001010;
            15'd28732: log10_cal = 16'b0000010111001010;
            15'd28733: log10_cal = 16'b0000010111001010;
            15'd28734: log10_cal = 16'b0000010111001010;
            15'd28735: log10_cal = 16'b0000010111001010;
            15'd28736: log10_cal = 16'b0000010111001010;
            15'd28737: log10_cal = 16'b0000010111001010;
            15'd28738: log10_cal = 16'b0000010111001010;
            15'd28739: log10_cal = 16'b0000010111001010;
            15'd28740: log10_cal = 16'b0000010111001010;
            15'd28741: log10_cal = 16'b0000010111001010;
            15'd28742: log10_cal = 16'b0000010111001010;
            15'd28743: log10_cal = 16'b0000010111001010;
            15'd28744: log10_cal = 16'b0000010111001011;
            15'd28745: log10_cal = 16'b0000010111001011;
            15'd28746: log10_cal = 16'b0000010111001011;
            15'd28747: log10_cal = 16'b0000010111001011;
            15'd28748: log10_cal = 16'b0000010111001011;
            15'd28749: log10_cal = 16'b0000010111001011;
            15'd28750: log10_cal = 16'b0000010111001011;
            15'd28751: log10_cal = 16'b0000010111001011;
            15'd28752: log10_cal = 16'b0000010111001011;
            15'd28753: log10_cal = 16'b0000010111001011;
            15'd28754: log10_cal = 16'b0000010111001011;
            15'd28755: log10_cal = 16'b0000010111001011;
            15'd28756: log10_cal = 16'b0000010111001011;
            15'd28757: log10_cal = 16'b0000010111001011;
            15'd28758: log10_cal = 16'b0000010111001011;
            15'd28759: log10_cal = 16'b0000010111001011;
            15'd28760: log10_cal = 16'b0000010111001011;
            15'd28761: log10_cal = 16'b0000010111001011;
            15'd28762: log10_cal = 16'b0000010111001011;
            15'd28763: log10_cal = 16'b0000010111001011;
            15'd28764: log10_cal = 16'b0000010111001011;
            15'd28765: log10_cal = 16'b0000010111001011;
            15'd28766: log10_cal = 16'b0000010111001011;
            15'd28767: log10_cal = 16'b0000010111001011;
            15'd28768: log10_cal = 16'b0000010111001011;
            15'd28769: log10_cal = 16'b0000010111001011;
            15'd28770: log10_cal = 16'b0000010111001011;
            15'd28771: log10_cal = 16'b0000010111001011;
            15'd28772: log10_cal = 16'b0000010111001011;
            15'd28773: log10_cal = 16'b0000010111001011;
            15'd28774: log10_cal = 16'b0000010111001011;
            15'd28775: log10_cal = 16'b0000010111001011;
            15'd28776: log10_cal = 16'b0000010111001011;
            15'd28777: log10_cal = 16'b0000010111001011;
            15'd28778: log10_cal = 16'b0000010111001011;
            15'd28779: log10_cal = 16'b0000010111001011;
            15'd28780: log10_cal = 16'b0000010111001011;
            15'd28781: log10_cal = 16'b0000010111001011;
            15'd28782: log10_cal = 16'b0000010111001011;
            15'd28783: log10_cal = 16'b0000010111001011;
            15'd28784: log10_cal = 16'b0000010111001011;
            15'd28785: log10_cal = 16'b0000010111001011;
            15'd28786: log10_cal = 16'b0000010111001011;
            15'd28787: log10_cal = 16'b0000010111001011;
            15'd28788: log10_cal = 16'b0000010111001011;
            15'd28789: log10_cal = 16'b0000010111001011;
            15'd28790: log10_cal = 16'b0000010111001011;
            15'd28791: log10_cal = 16'b0000010111001011;
            15'd28792: log10_cal = 16'b0000010111001011;
            15'd28793: log10_cal = 16'b0000010111001011;
            15'd28794: log10_cal = 16'b0000010111001011;
            15'd28795: log10_cal = 16'b0000010111001011;
            15'd28796: log10_cal = 16'b0000010111001011;
            15'd28797: log10_cal = 16'b0000010111001011;
            15'd28798: log10_cal = 16'b0000010111001011;
            15'd28799: log10_cal = 16'b0000010111001011;
            15'd28800: log10_cal = 16'b0000010111001011;
            15'd28801: log10_cal = 16'b0000010111001011;
            15'd28802: log10_cal = 16'b0000010111001011;
            15'd28803: log10_cal = 16'b0000010111001011;
            15'd28804: log10_cal = 16'b0000010111001011;
            15'd28805: log10_cal = 16'b0000010111001011;
            15'd28806: log10_cal = 16'b0000010111001011;
            15'd28807: log10_cal = 16'b0000010111001011;
            15'd28808: log10_cal = 16'b0000010111001011;
            15'd28809: log10_cal = 16'b0000010111001100;
            15'd28810: log10_cal = 16'b0000010111001100;
            15'd28811: log10_cal = 16'b0000010111001100;
            15'd28812: log10_cal = 16'b0000010111001100;
            15'd28813: log10_cal = 16'b0000010111001100;
            15'd28814: log10_cal = 16'b0000010111001100;
            15'd28815: log10_cal = 16'b0000010111001100;
            15'd28816: log10_cal = 16'b0000010111001100;
            15'd28817: log10_cal = 16'b0000010111001100;
            15'd28818: log10_cal = 16'b0000010111001100;
            15'd28819: log10_cal = 16'b0000010111001100;
            15'd28820: log10_cal = 16'b0000010111001100;
            15'd28821: log10_cal = 16'b0000010111001100;
            15'd28822: log10_cal = 16'b0000010111001100;
            15'd28823: log10_cal = 16'b0000010111001100;
            15'd28824: log10_cal = 16'b0000010111001100;
            15'd28825: log10_cal = 16'b0000010111001100;
            15'd28826: log10_cal = 16'b0000010111001100;
            15'd28827: log10_cal = 16'b0000010111001100;
            15'd28828: log10_cal = 16'b0000010111001100;
            15'd28829: log10_cal = 16'b0000010111001100;
            15'd28830: log10_cal = 16'b0000010111001100;
            15'd28831: log10_cal = 16'b0000010111001100;
            15'd28832: log10_cal = 16'b0000010111001100;
            15'd28833: log10_cal = 16'b0000010111001100;
            15'd28834: log10_cal = 16'b0000010111001100;
            15'd28835: log10_cal = 16'b0000010111001100;
            15'd28836: log10_cal = 16'b0000010111001100;
            15'd28837: log10_cal = 16'b0000010111001100;
            15'd28838: log10_cal = 16'b0000010111001100;
            15'd28839: log10_cal = 16'b0000010111001100;
            15'd28840: log10_cal = 16'b0000010111001100;
            15'd28841: log10_cal = 16'b0000010111001100;
            15'd28842: log10_cal = 16'b0000010111001100;
            15'd28843: log10_cal = 16'b0000010111001100;
            15'd28844: log10_cal = 16'b0000010111001100;
            15'd28845: log10_cal = 16'b0000010111001100;
            15'd28846: log10_cal = 16'b0000010111001100;
            15'd28847: log10_cal = 16'b0000010111001100;
            15'd28848: log10_cal = 16'b0000010111001100;
            15'd28849: log10_cal = 16'b0000010111001100;
            15'd28850: log10_cal = 16'b0000010111001100;
            15'd28851: log10_cal = 16'b0000010111001100;
            15'd28852: log10_cal = 16'b0000010111001100;
            15'd28853: log10_cal = 16'b0000010111001100;
            15'd28854: log10_cal = 16'b0000010111001100;
            15'd28855: log10_cal = 16'b0000010111001100;
            15'd28856: log10_cal = 16'b0000010111001100;
            15'd28857: log10_cal = 16'b0000010111001100;
            15'd28858: log10_cal = 16'b0000010111001100;
            15'd28859: log10_cal = 16'b0000010111001100;
            15'd28860: log10_cal = 16'b0000010111001100;
            15'd28861: log10_cal = 16'b0000010111001100;
            15'd28862: log10_cal = 16'b0000010111001100;
            15'd28863: log10_cal = 16'b0000010111001100;
            15'd28864: log10_cal = 16'b0000010111001100;
            15'd28865: log10_cal = 16'b0000010111001100;
            15'd28866: log10_cal = 16'b0000010111001100;
            15'd28867: log10_cal = 16'b0000010111001100;
            15'd28868: log10_cal = 16'b0000010111001100;
            15'd28869: log10_cal = 16'b0000010111001100;
            15'd28870: log10_cal = 16'b0000010111001100;
            15'd28871: log10_cal = 16'b0000010111001100;
            15'd28872: log10_cal = 16'b0000010111001100;
            15'd28873: log10_cal = 16'b0000010111001100;
            15'd28874: log10_cal = 16'b0000010111001101;
            15'd28875: log10_cal = 16'b0000010111001101;
            15'd28876: log10_cal = 16'b0000010111001101;
            15'd28877: log10_cal = 16'b0000010111001101;
            15'd28878: log10_cal = 16'b0000010111001101;
            15'd28879: log10_cal = 16'b0000010111001101;
            15'd28880: log10_cal = 16'b0000010111001101;
            15'd28881: log10_cal = 16'b0000010111001101;
            15'd28882: log10_cal = 16'b0000010111001101;
            15'd28883: log10_cal = 16'b0000010111001101;
            15'd28884: log10_cal = 16'b0000010111001101;
            15'd28885: log10_cal = 16'b0000010111001101;
            15'd28886: log10_cal = 16'b0000010111001101;
            15'd28887: log10_cal = 16'b0000010111001101;
            15'd28888: log10_cal = 16'b0000010111001101;
            15'd28889: log10_cal = 16'b0000010111001101;
            15'd28890: log10_cal = 16'b0000010111001101;
            15'd28891: log10_cal = 16'b0000010111001101;
            15'd28892: log10_cal = 16'b0000010111001101;
            15'd28893: log10_cal = 16'b0000010111001101;
            15'd28894: log10_cal = 16'b0000010111001101;
            15'd28895: log10_cal = 16'b0000010111001101;
            15'd28896: log10_cal = 16'b0000010111001101;
            15'd28897: log10_cal = 16'b0000010111001101;
            15'd28898: log10_cal = 16'b0000010111001101;
            15'd28899: log10_cal = 16'b0000010111001101;
            15'd28900: log10_cal = 16'b0000010111001101;
            15'd28901: log10_cal = 16'b0000010111001101;
            15'd28902: log10_cal = 16'b0000010111001101;
            15'd28903: log10_cal = 16'b0000010111001101;
            15'd28904: log10_cal = 16'b0000010111001101;
            15'd28905: log10_cal = 16'b0000010111001101;
            15'd28906: log10_cal = 16'b0000010111001101;
            15'd28907: log10_cal = 16'b0000010111001101;
            15'd28908: log10_cal = 16'b0000010111001101;
            15'd28909: log10_cal = 16'b0000010111001101;
            15'd28910: log10_cal = 16'b0000010111001101;
            15'd28911: log10_cal = 16'b0000010111001101;
            15'd28912: log10_cal = 16'b0000010111001101;
            15'd28913: log10_cal = 16'b0000010111001101;
            15'd28914: log10_cal = 16'b0000010111001101;
            15'd28915: log10_cal = 16'b0000010111001101;
            15'd28916: log10_cal = 16'b0000010111001101;
            15'd28917: log10_cal = 16'b0000010111001101;
            15'd28918: log10_cal = 16'b0000010111001101;
            15'd28919: log10_cal = 16'b0000010111001101;
            15'd28920: log10_cal = 16'b0000010111001101;
            15'd28921: log10_cal = 16'b0000010111001101;
            15'd28922: log10_cal = 16'b0000010111001101;
            15'd28923: log10_cal = 16'b0000010111001101;
            15'd28924: log10_cal = 16'b0000010111001101;
            15'd28925: log10_cal = 16'b0000010111001101;
            15'd28926: log10_cal = 16'b0000010111001101;
            15'd28927: log10_cal = 16'b0000010111001101;
            15'd28928: log10_cal = 16'b0000010111001101;
            15'd28929: log10_cal = 16'b0000010111001101;
            15'd28930: log10_cal = 16'b0000010111001101;
            15'd28931: log10_cal = 16'b0000010111001101;
            15'd28932: log10_cal = 16'b0000010111001101;
            15'd28933: log10_cal = 16'b0000010111001101;
            15'd28934: log10_cal = 16'b0000010111001101;
            15'd28935: log10_cal = 16'b0000010111001101;
            15'd28936: log10_cal = 16'b0000010111001101;
            15'd28937: log10_cal = 16'b0000010111001101;
            15'd28938: log10_cal = 16'b0000010111001101;
            15'd28939: log10_cal = 16'b0000010111001110;
            15'd28940: log10_cal = 16'b0000010111001110;
            15'd28941: log10_cal = 16'b0000010111001110;
            15'd28942: log10_cal = 16'b0000010111001110;
            15'd28943: log10_cal = 16'b0000010111001110;
            15'd28944: log10_cal = 16'b0000010111001110;
            15'd28945: log10_cal = 16'b0000010111001110;
            15'd28946: log10_cal = 16'b0000010111001110;
            15'd28947: log10_cal = 16'b0000010111001110;
            15'd28948: log10_cal = 16'b0000010111001110;
            15'd28949: log10_cal = 16'b0000010111001110;
            15'd28950: log10_cal = 16'b0000010111001110;
            15'd28951: log10_cal = 16'b0000010111001110;
            15'd28952: log10_cal = 16'b0000010111001110;
            15'd28953: log10_cal = 16'b0000010111001110;
            15'd28954: log10_cal = 16'b0000010111001110;
            15'd28955: log10_cal = 16'b0000010111001110;
            15'd28956: log10_cal = 16'b0000010111001110;
            15'd28957: log10_cal = 16'b0000010111001110;
            15'd28958: log10_cal = 16'b0000010111001110;
            15'd28959: log10_cal = 16'b0000010111001110;
            15'd28960: log10_cal = 16'b0000010111001110;
            15'd28961: log10_cal = 16'b0000010111001110;
            15'd28962: log10_cal = 16'b0000010111001110;
            15'd28963: log10_cal = 16'b0000010111001110;
            15'd28964: log10_cal = 16'b0000010111001110;
            15'd28965: log10_cal = 16'b0000010111001110;
            15'd28966: log10_cal = 16'b0000010111001110;
            15'd28967: log10_cal = 16'b0000010111001110;
            15'd28968: log10_cal = 16'b0000010111001110;
            15'd28969: log10_cal = 16'b0000010111001110;
            15'd28970: log10_cal = 16'b0000010111001110;
            15'd28971: log10_cal = 16'b0000010111001110;
            15'd28972: log10_cal = 16'b0000010111001110;
            15'd28973: log10_cal = 16'b0000010111001110;
            15'd28974: log10_cal = 16'b0000010111001110;
            15'd28975: log10_cal = 16'b0000010111001110;
            15'd28976: log10_cal = 16'b0000010111001110;
            15'd28977: log10_cal = 16'b0000010111001110;
            15'd28978: log10_cal = 16'b0000010111001110;
            15'd28979: log10_cal = 16'b0000010111001110;
            15'd28980: log10_cal = 16'b0000010111001110;
            15'd28981: log10_cal = 16'b0000010111001110;
            15'd28982: log10_cal = 16'b0000010111001110;
            15'd28983: log10_cal = 16'b0000010111001110;
            15'd28984: log10_cal = 16'b0000010111001110;
            15'd28985: log10_cal = 16'b0000010111001110;
            15'd28986: log10_cal = 16'b0000010111001110;
            15'd28987: log10_cal = 16'b0000010111001110;
            15'd28988: log10_cal = 16'b0000010111001110;
            15'd28989: log10_cal = 16'b0000010111001110;
            15'd28990: log10_cal = 16'b0000010111001110;
            15'd28991: log10_cal = 16'b0000010111001110;
            15'd28992: log10_cal = 16'b0000010111001110;
            15'd28993: log10_cal = 16'b0000010111001110;
            15'd28994: log10_cal = 16'b0000010111001110;
            15'd28995: log10_cal = 16'b0000010111001110;
            15'd28996: log10_cal = 16'b0000010111001110;
            15'd28997: log10_cal = 16'b0000010111001110;
            15'd28998: log10_cal = 16'b0000010111001110;
            15'd28999: log10_cal = 16'b0000010111001110;
            15'd29000: log10_cal = 16'b0000010111001110;
            15'd29001: log10_cal = 16'b0000010111001110;
            15'd29002: log10_cal = 16'b0000010111001110;
            15'd29003: log10_cal = 16'b0000010111001110;
            15'd29004: log10_cal = 16'b0000010111001111;
            15'd29005: log10_cal = 16'b0000010111001111;
            15'd29006: log10_cal = 16'b0000010111001111;
            15'd29007: log10_cal = 16'b0000010111001111;
            15'd29008: log10_cal = 16'b0000010111001111;
            15'd29009: log10_cal = 16'b0000010111001111;
            15'd29010: log10_cal = 16'b0000010111001111;
            15'd29011: log10_cal = 16'b0000010111001111;
            15'd29012: log10_cal = 16'b0000010111001111;
            15'd29013: log10_cal = 16'b0000010111001111;
            15'd29014: log10_cal = 16'b0000010111001111;
            15'd29015: log10_cal = 16'b0000010111001111;
            15'd29016: log10_cal = 16'b0000010111001111;
            15'd29017: log10_cal = 16'b0000010111001111;
            15'd29018: log10_cal = 16'b0000010111001111;
            15'd29019: log10_cal = 16'b0000010111001111;
            15'd29020: log10_cal = 16'b0000010111001111;
            15'd29021: log10_cal = 16'b0000010111001111;
            15'd29022: log10_cal = 16'b0000010111001111;
            15'd29023: log10_cal = 16'b0000010111001111;
            15'd29024: log10_cal = 16'b0000010111001111;
            15'd29025: log10_cal = 16'b0000010111001111;
            15'd29026: log10_cal = 16'b0000010111001111;
            15'd29027: log10_cal = 16'b0000010111001111;
            15'd29028: log10_cal = 16'b0000010111001111;
            15'd29029: log10_cal = 16'b0000010111001111;
            15'd29030: log10_cal = 16'b0000010111001111;
            15'd29031: log10_cal = 16'b0000010111001111;
            15'd29032: log10_cal = 16'b0000010111001111;
            15'd29033: log10_cal = 16'b0000010111001111;
            15'd29034: log10_cal = 16'b0000010111001111;
            15'd29035: log10_cal = 16'b0000010111001111;
            15'd29036: log10_cal = 16'b0000010111001111;
            15'd29037: log10_cal = 16'b0000010111001111;
            15'd29038: log10_cal = 16'b0000010111001111;
            15'd29039: log10_cal = 16'b0000010111001111;
            15'd29040: log10_cal = 16'b0000010111001111;
            15'd29041: log10_cal = 16'b0000010111001111;
            15'd29042: log10_cal = 16'b0000010111001111;
            15'd29043: log10_cal = 16'b0000010111001111;
            15'd29044: log10_cal = 16'b0000010111001111;
            15'd29045: log10_cal = 16'b0000010111001111;
            15'd29046: log10_cal = 16'b0000010111001111;
            15'd29047: log10_cal = 16'b0000010111001111;
            15'd29048: log10_cal = 16'b0000010111001111;
            15'd29049: log10_cal = 16'b0000010111001111;
            15'd29050: log10_cal = 16'b0000010111001111;
            15'd29051: log10_cal = 16'b0000010111001111;
            15'd29052: log10_cal = 16'b0000010111001111;
            15'd29053: log10_cal = 16'b0000010111001111;
            15'd29054: log10_cal = 16'b0000010111001111;
            15'd29055: log10_cal = 16'b0000010111001111;
            15'd29056: log10_cal = 16'b0000010111001111;
            15'd29057: log10_cal = 16'b0000010111001111;
            15'd29058: log10_cal = 16'b0000010111001111;
            15'd29059: log10_cal = 16'b0000010111001111;
            15'd29060: log10_cal = 16'b0000010111001111;
            15'd29061: log10_cal = 16'b0000010111001111;
            15'd29062: log10_cal = 16'b0000010111001111;
            15'd29063: log10_cal = 16'b0000010111001111;
            15'd29064: log10_cal = 16'b0000010111001111;
            15'd29065: log10_cal = 16'b0000010111001111;
            15'd29066: log10_cal = 16'b0000010111001111;
            15'd29067: log10_cal = 16'b0000010111001111;
            15'd29068: log10_cal = 16'b0000010111001111;
            15'd29069: log10_cal = 16'b0000010111010000;
            15'd29070: log10_cal = 16'b0000010111010000;
            15'd29071: log10_cal = 16'b0000010111010000;
            15'd29072: log10_cal = 16'b0000010111010000;
            15'd29073: log10_cal = 16'b0000010111010000;
            15'd29074: log10_cal = 16'b0000010111010000;
            15'd29075: log10_cal = 16'b0000010111010000;
            15'd29076: log10_cal = 16'b0000010111010000;
            15'd29077: log10_cal = 16'b0000010111010000;
            15'd29078: log10_cal = 16'b0000010111010000;
            15'd29079: log10_cal = 16'b0000010111010000;
            15'd29080: log10_cal = 16'b0000010111010000;
            15'd29081: log10_cal = 16'b0000010111010000;
            15'd29082: log10_cal = 16'b0000010111010000;
            15'd29083: log10_cal = 16'b0000010111010000;
            15'd29084: log10_cal = 16'b0000010111010000;
            15'd29085: log10_cal = 16'b0000010111010000;
            15'd29086: log10_cal = 16'b0000010111010000;
            15'd29087: log10_cal = 16'b0000010111010000;
            15'd29088: log10_cal = 16'b0000010111010000;
            15'd29089: log10_cal = 16'b0000010111010000;
            15'd29090: log10_cal = 16'b0000010111010000;
            15'd29091: log10_cal = 16'b0000010111010000;
            15'd29092: log10_cal = 16'b0000010111010000;
            15'd29093: log10_cal = 16'b0000010111010000;
            15'd29094: log10_cal = 16'b0000010111010000;
            15'd29095: log10_cal = 16'b0000010111010000;
            15'd29096: log10_cal = 16'b0000010111010000;
            15'd29097: log10_cal = 16'b0000010111010000;
            15'd29098: log10_cal = 16'b0000010111010000;
            15'd29099: log10_cal = 16'b0000010111010000;
            15'd29100: log10_cal = 16'b0000010111010000;
            15'd29101: log10_cal = 16'b0000010111010000;
            15'd29102: log10_cal = 16'b0000010111010000;
            15'd29103: log10_cal = 16'b0000010111010000;
            15'd29104: log10_cal = 16'b0000010111010000;
            15'd29105: log10_cal = 16'b0000010111010000;
            15'd29106: log10_cal = 16'b0000010111010000;
            15'd29107: log10_cal = 16'b0000010111010000;
            15'd29108: log10_cal = 16'b0000010111010000;
            15'd29109: log10_cal = 16'b0000010111010000;
            15'd29110: log10_cal = 16'b0000010111010000;
            15'd29111: log10_cal = 16'b0000010111010000;
            15'd29112: log10_cal = 16'b0000010111010000;
            15'd29113: log10_cal = 16'b0000010111010000;
            15'd29114: log10_cal = 16'b0000010111010000;
            15'd29115: log10_cal = 16'b0000010111010000;
            15'd29116: log10_cal = 16'b0000010111010000;
            15'd29117: log10_cal = 16'b0000010111010000;
            15'd29118: log10_cal = 16'b0000010111010000;
            15'd29119: log10_cal = 16'b0000010111010000;
            15'd29120: log10_cal = 16'b0000010111010000;
            15'd29121: log10_cal = 16'b0000010111010000;
            15'd29122: log10_cal = 16'b0000010111010000;
            15'd29123: log10_cal = 16'b0000010111010000;
            15'd29124: log10_cal = 16'b0000010111010000;
            15'd29125: log10_cal = 16'b0000010111010000;
            15'd29126: log10_cal = 16'b0000010111010000;
            15'd29127: log10_cal = 16'b0000010111010000;
            15'd29128: log10_cal = 16'b0000010111010000;
            15'd29129: log10_cal = 16'b0000010111010000;
            15'd29130: log10_cal = 16'b0000010111010000;
            15'd29131: log10_cal = 16'b0000010111010000;
            15'd29132: log10_cal = 16'b0000010111010000;
            15'd29133: log10_cal = 16'b0000010111010000;
            15'd29134: log10_cal = 16'b0000010111010000;
            15'd29135: log10_cal = 16'b0000010111010001;
            15'd29136: log10_cal = 16'b0000010111010001;
            15'd29137: log10_cal = 16'b0000010111010001;
            15'd29138: log10_cal = 16'b0000010111010001;
            15'd29139: log10_cal = 16'b0000010111010001;
            15'd29140: log10_cal = 16'b0000010111010001;
            15'd29141: log10_cal = 16'b0000010111010001;
            15'd29142: log10_cal = 16'b0000010111010001;
            15'd29143: log10_cal = 16'b0000010111010001;
            15'd29144: log10_cal = 16'b0000010111010001;
            15'd29145: log10_cal = 16'b0000010111010001;
            15'd29146: log10_cal = 16'b0000010111010001;
            15'd29147: log10_cal = 16'b0000010111010001;
            15'd29148: log10_cal = 16'b0000010111010001;
            15'd29149: log10_cal = 16'b0000010111010001;
            15'd29150: log10_cal = 16'b0000010111010001;
            15'd29151: log10_cal = 16'b0000010111010001;
            15'd29152: log10_cal = 16'b0000010111010001;
            15'd29153: log10_cal = 16'b0000010111010001;
            15'd29154: log10_cal = 16'b0000010111010001;
            15'd29155: log10_cal = 16'b0000010111010001;
            15'd29156: log10_cal = 16'b0000010111010001;
            15'd29157: log10_cal = 16'b0000010111010001;
            15'd29158: log10_cal = 16'b0000010111010001;
            15'd29159: log10_cal = 16'b0000010111010001;
            15'd29160: log10_cal = 16'b0000010111010001;
            15'd29161: log10_cal = 16'b0000010111010001;
            15'd29162: log10_cal = 16'b0000010111010001;
            15'd29163: log10_cal = 16'b0000010111010001;
            15'd29164: log10_cal = 16'b0000010111010001;
            15'd29165: log10_cal = 16'b0000010111010001;
            15'd29166: log10_cal = 16'b0000010111010001;
            15'd29167: log10_cal = 16'b0000010111010001;
            15'd29168: log10_cal = 16'b0000010111010001;
            15'd29169: log10_cal = 16'b0000010111010001;
            15'd29170: log10_cal = 16'b0000010111010001;
            15'd29171: log10_cal = 16'b0000010111010001;
            15'd29172: log10_cal = 16'b0000010111010001;
            15'd29173: log10_cal = 16'b0000010111010001;
            15'd29174: log10_cal = 16'b0000010111010001;
            15'd29175: log10_cal = 16'b0000010111010001;
            15'd29176: log10_cal = 16'b0000010111010001;
            15'd29177: log10_cal = 16'b0000010111010001;
            15'd29178: log10_cal = 16'b0000010111010001;
            15'd29179: log10_cal = 16'b0000010111010001;
            15'd29180: log10_cal = 16'b0000010111010001;
            15'd29181: log10_cal = 16'b0000010111010001;
            15'd29182: log10_cal = 16'b0000010111010001;
            15'd29183: log10_cal = 16'b0000010111010001;
            15'd29184: log10_cal = 16'b0000010111010001;
            15'd29185: log10_cal = 16'b0000010111010001;
            15'd29186: log10_cal = 16'b0000010111010001;
            15'd29187: log10_cal = 16'b0000010111010001;
            15'd29188: log10_cal = 16'b0000010111010001;
            15'd29189: log10_cal = 16'b0000010111010001;
            15'd29190: log10_cal = 16'b0000010111010001;
            15'd29191: log10_cal = 16'b0000010111010001;
            15'd29192: log10_cal = 16'b0000010111010001;
            15'd29193: log10_cal = 16'b0000010111010001;
            15'd29194: log10_cal = 16'b0000010111010001;
            15'd29195: log10_cal = 16'b0000010111010001;
            15'd29196: log10_cal = 16'b0000010111010001;
            15'd29197: log10_cal = 16'b0000010111010001;
            15'd29198: log10_cal = 16'b0000010111010001;
            15'd29199: log10_cal = 16'b0000010111010001;
            15'd29200: log10_cal = 16'b0000010111010010;
            15'd29201: log10_cal = 16'b0000010111010010;
            15'd29202: log10_cal = 16'b0000010111010010;
            15'd29203: log10_cal = 16'b0000010111010010;
            15'd29204: log10_cal = 16'b0000010111010010;
            15'd29205: log10_cal = 16'b0000010111010010;
            15'd29206: log10_cal = 16'b0000010111010010;
            15'd29207: log10_cal = 16'b0000010111010010;
            15'd29208: log10_cal = 16'b0000010111010010;
            15'd29209: log10_cal = 16'b0000010111010010;
            15'd29210: log10_cal = 16'b0000010111010010;
            15'd29211: log10_cal = 16'b0000010111010010;
            15'd29212: log10_cal = 16'b0000010111010010;
            15'd29213: log10_cal = 16'b0000010111010010;
            15'd29214: log10_cal = 16'b0000010111010010;
            15'd29215: log10_cal = 16'b0000010111010010;
            15'd29216: log10_cal = 16'b0000010111010010;
            15'd29217: log10_cal = 16'b0000010111010010;
            15'd29218: log10_cal = 16'b0000010111010010;
            15'd29219: log10_cal = 16'b0000010111010010;
            15'd29220: log10_cal = 16'b0000010111010010;
            15'd29221: log10_cal = 16'b0000010111010010;
            15'd29222: log10_cal = 16'b0000010111010010;
            15'd29223: log10_cal = 16'b0000010111010010;
            15'd29224: log10_cal = 16'b0000010111010010;
            15'd29225: log10_cal = 16'b0000010111010010;
            15'd29226: log10_cal = 16'b0000010111010010;
            15'd29227: log10_cal = 16'b0000010111010010;
            15'd29228: log10_cal = 16'b0000010111010010;
            15'd29229: log10_cal = 16'b0000010111010010;
            15'd29230: log10_cal = 16'b0000010111010010;
            15'd29231: log10_cal = 16'b0000010111010010;
            15'd29232: log10_cal = 16'b0000010111010010;
            15'd29233: log10_cal = 16'b0000010111010010;
            15'd29234: log10_cal = 16'b0000010111010010;
            15'd29235: log10_cal = 16'b0000010111010010;
            15'd29236: log10_cal = 16'b0000010111010010;
            15'd29237: log10_cal = 16'b0000010111010010;
            15'd29238: log10_cal = 16'b0000010111010010;
            15'd29239: log10_cal = 16'b0000010111010010;
            15'd29240: log10_cal = 16'b0000010111010010;
            15'd29241: log10_cal = 16'b0000010111010010;
            15'd29242: log10_cal = 16'b0000010111010010;
            15'd29243: log10_cal = 16'b0000010111010010;
            15'd29244: log10_cal = 16'b0000010111010010;
            15'd29245: log10_cal = 16'b0000010111010010;
            15'd29246: log10_cal = 16'b0000010111010010;
            15'd29247: log10_cal = 16'b0000010111010010;
            15'd29248: log10_cal = 16'b0000010111010010;
            15'd29249: log10_cal = 16'b0000010111010010;
            15'd29250: log10_cal = 16'b0000010111010010;
            15'd29251: log10_cal = 16'b0000010111010010;
            15'd29252: log10_cal = 16'b0000010111010010;
            15'd29253: log10_cal = 16'b0000010111010010;
            15'd29254: log10_cal = 16'b0000010111010010;
            15'd29255: log10_cal = 16'b0000010111010010;
            15'd29256: log10_cal = 16'b0000010111010010;
            15'd29257: log10_cal = 16'b0000010111010010;
            15'd29258: log10_cal = 16'b0000010111010010;
            15'd29259: log10_cal = 16'b0000010111010010;
            15'd29260: log10_cal = 16'b0000010111010010;
            15'd29261: log10_cal = 16'b0000010111010010;
            15'd29262: log10_cal = 16'b0000010111010010;
            15'd29263: log10_cal = 16'b0000010111010010;
            15'd29264: log10_cal = 16'b0000010111010010;
            15'd29265: log10_cal = 16'b0000010111010010;
            15'd29266: log10_cal = 16'b0000010111010011;
            15'd29267: log10_cal = 16'b0000010111010011;
            15'd29268: log10_cal = 16'b0000010111010011;
            15'd29269: log10_cal = 16'b0000010111010011;
            15'd29270: log10_cal = 16'b0000010111010011;
            15'd29271: log10_cal = 16'b0000010111010011;
            15'd29272: log10_cal = 16'b0000010111010011;
            15'd29273: log10_cal = 16'b0000010111010011;
            15'd29274: log10_cal = 16'b0000010111010011;
            15'd29275: log10_cal = 16'b0000010111010011;
            15'd29276: log10_cal = 16'b0000010111010011;
            15'd29277: log10_cal = 16'b0000010111010011;
            15'd29278: log10_cal = 16'b0000010111010011;
            15'd29279: log10_cal = 16'b0000010111010011;
            15'd29280: log10_cal = 16'b0000010111010011;
            15'd29281: log10_cal = 16'b0000010111010011;
            15'd29282: log10_cal = 16'b0000010111010011;
            15'd29283: log10_cal = 16'b0000010111010011;
            15'd29284: log10_cal = 16'b0000010111010011;
            15'd29285: log10_cal = 16'b0000010111010011;
            15'd29286: log10_cal = 16'b0000010111010011;
            15'd29287: log10_cal = 16'b0000010111010011;
            15'd29288: log10_cal = 16'b0000010111010011;
            15'd29289: log10_cal = 16'b0000010111010011;
            15'd29290: log10_cal = 16'b0000010111010011;
            15'd29291: log10_cal = 16'b0000010111010011;
            15'd29292: log10_cal = 16'b0000010111010011;
            15'd29293: log10_cal = 16'b0000010111010011;
            15'd29294: log10_cal = 16'b0000010111010011;
            15'd29295: log10_cal = 16'b0000010111010011;
            15'd29296: log10_cal = 16'b0000010111010011;
            15'd29297: log10_cal = 16'b0000010111010011;
            15'd29298: log10_cal = 16'b0000010111010011;
            15'd29299: log10_cal = 16'b0000010111010011;
            15'd29300: log10_cal = 16'b0000010111010011;
            15'd29301: log10_cal = 16'b0000010111010011;
            15'd29302: log10_cal = 16'b0000010111010011;
            15'd29303: log10_cal = 16'b0000010111010011;
            15'd29304: log10_cal = 16'b0000010111010011;
            15'd29305: log10_cal = 16'b0000010111010011;
            15'd29306: log10_cal = 16'b0000010111010011;
            15'd29307: log10_cal = 16'b0000010111010011;
            15'd29308: log10_cal = 16'b0000010111010011;
            15'd29309: log10_cal = 16'b0000010111010011;
            15'd29310: log10_cal = 16'b0000010111010011;
            15'd29311: log10_cal = 16'b0000010111010011;
            15'd29312: log10_cal = 16'b0000010111010011;
            15'd29313: log10_cal = 16'b0000010111010011;
            15'd29314: log10_cal = 16'b0000010111010011;
            15'd29315: log10_cal = 16'b0000010111010011;
            15'd29316: log10_cal = 16'b0000010111010011;
            15'd29317: log10_cal = 16'b0000010111010011;
            15'd29318: log10_cal = 16'b0000010111010011;
            15'd29319: log10_cal = 16'b0000010111010011;
            15'd29320: log10_cal = 16'b0000010111010011;
            15'd29321: log10_cal = 16'b0000010111010011;
            15'd29322: log10_cal = 16'b0000010111010011;
            15'd29323: log10_cal = 16'b0000010111010011;
            15'd29324: log10_cal = 16'b0000010111010011;
            15'd29325: log10_cal = 16'b0000010111010011;
            15'd29326: log10_cal = 16'b0000010111010011;
            15'd29327: log10_cal = 16'b0000010111010011;
            15'd29328: log10_cal = 16'b0000010111010011;
            15'd29329: log10_cal = 16'b0000010111010011;
            15'd29330: log10_cal = 16'b0000010111010011;
            15'd29331: log10_cal = 16'b0000010111010011;
            15'd29332: log10_cal = 16'b0000010111010100;
            15'd29333: log10_cal = 16'b0000010111010100;
            15'd29334: log10_cal = 16'b0000010111010100;
            15'd29335: log10_cal = 16'b0000010111010100;
            15'd29336: log10_cal = 16'b0000010111010100;
            15'd29337: log10_cal = 16'b0000010111010100;
            15'd29338: log10_cal = 16'b0000010111010100;
            15'd29339: log10_cal = 16'b0000010111010100;
            15'd29340: log10_cal = 16'b0000010111010100;
            15'd29341: log10_cal = 16'b0000010111010100;
            15'd29342: log10_cal = 16'b0000010111010100;
            15'd29343: log10_cal = 16'b0000010111010100;
            15'd29344: log10_cal = 16'b0000010111010100;
            15'd29345: log10_cal = 16'b0000010111010100;
            15'd29346: log10_cal = 16'b0000010111010100;
            15'd29347: log10_cal = 16'b0000010111010100;
            15'd29348: log10_cal = 16'b0000010111010100;
            15'd29349: log10_cal = 16'b0000010111010100;
            15'd29350: log10_cal = 16'b0000010111010100;
            15'd29351: log10_cal = 16'b0000010111010100;
            15'd29352: log10_cal = 16'b0000010111010100;
            15'd29353: log10_cal = 16'b0000010111010100;
            15'd29354: log10_cal = 16'b0000010111010100;
            15'd29355: log10_cal = 16'b0000010111010100;
            15'd29356: log10_cal = 16'b0000010111010100;
            15'd29357: log10_cal = 16'b0000010111010100;
            15'd29358: log10_cal = 16'b0000010111010100;
            15'd29359: log10_cal = 16'b0000010111010100;
            15'd29360: log10_cal = 16'b0000010111010100;
            15'd29361: log10_cal = 16'b0000010111010100;
            15'd29362: log10_cal = 16'b0000010111010100;
            15'd29363: log10_cal = 16'b0000010111010100;
            15'd29364: log10_cal = 16'b0000010111010100;
            15'd29365: log10_cal = 16'b0000010111010100;
            15'd29366: log10_cal = 16'b0000010111010100;
            15'd29367: log10_cal = 16'b0000010111010100;
            15'd29368: log10_cal = 16'b0000010111010100;
            15'd29369: log10_cal = 16'b0000010111010100;
            15'd29370: log10_cal = 16'b0000010111010100;
            15'd29371: log10_cal = 16'b0000010111010100;
            15'd29372: log10_cal = 16'b0000010111010100;
            15'd29373: log10_cal = 16'b0000010111010100;
            15'd29374: log10_cal = 16'b0000010111010100;
            15'd29375: log10_cal = 16'b0000010111010100;
            15'd29376: log10_cal = 16'b0000010111010100;
            15'd29377: log10_cal = 16'b0000010111010100;
            15'd29378: log10_cal = 16'b0000010111010100;
            15'd29379: log10_cal = 16'b0000010111010100;
            15'd29380: log10_cal = 16'b0000010111010100;
            15'd29381: log10_cal = 16'b0000010111010100;
            15'd29382: log10_cal = 16'b0000010111010100;
            15'd29383: log10_cal = 16'b0000010111010100;
            15'd29384: log10_cal = 16'b0000010111010100;
            15'd29385: log10_cal = 16'b0000010111010100;
            15'd29386: log10_cal = 16'b0000010111010100;
            15'd29387: log10_cal = 16'b0000010111010100;
            15'd29388: log10_cal = 16'b0000010111010100;
            15'd29389: log10_cal = 16'b0000010111010100;
            15'd29390: log10_cal = 16'b0000010111010100;
            15'd29391: log10_cal = 16'b0000010111010100;
            15'd29392: log10_cal = 16'b0000010111010100;
            15'd29393: log10_cal = 16'b0000010111010100;
            15'd29394: log10_cal = 16'b0000010111010100;
            15'd29395: log10_cal = 16'b0000010111010100;
            15'd29396: log10_cal = 16'b0000010111010100;
            15'd29397: log10_cal = 16'b0000010111010100;
            15'd29398: log10_cal = 16'b0000010111010101;
            15'd29399: log10_cal = 16'b0000010111010101;
            15'd29400: log10_cal = 16'b0000010111010101;
            15'd29401: log10_cal = 16'b0000010111010101;
            15'd29402: log10_cal = 16'b0000010111010101;
            15'd29403: log10_cal = 16'b0000010111010101;
            15'd29404: log10_cal = 16'b0000010111010101;
            15'd29405: log10_cal = 16'b0000010111010101;
            15'd29406: log10_cal = 16'b0000010111010101;
            15'd29407: log10_cal = 16'b0000010111010101;
            15'd29408: log10_cal = 16'b0000010111010101;
            15'd29409: log10_cal = 16'b0000010111010101;
            15'd29410: log10_cal = 16'b0000010111010101;
            15'd29411: log10_cal = 16'b0000010111010101;
            15'd29412: log10_cal = 16'b0000010111010101;
            15'd29413: log10_cal = 16'b0000010111010101;
            15'd29414: log10_cal = 16'b0000010111010101;
            15'd29415: log10_cal = 16'b0000010111010101;
            15'd29416: log10_cal = 16'b0000010111010101;
            15'd29417: log10_cal = 16'b0000010111010101;
            15'd29418: log10_cal = 16'b0000010111010101;
            15'd29419: log10_cal = 16'b0000010111010101;
            15'd29420: log10_cal = 16'b0000010111010101;
            15'd29421: log10_cal = 16'b0000010111010101;
            15'd29422: log10_cal = 16'b0000010111010101;
            15'd29423: log10_cal = 16'b0000010111010101;
            15'd29424: log10_cal = 16'b0000010111010101;
            15'd29425: log10_cal = 16'b0000010111010101;
            15'd29426: log10_cal = 16'b0000010111010101;
            15'd29427: log10_cal = 16'b0000010111010101;
            15'd29428: log10_cal = 16'b0000010111010101;
            15'd29429: log10_cal = 16'b0000010111010101;
            15'd29430: log10_cal = 16'b0000010111010101;
            15'd29431: log10_cal = 16'b0000010111010101;
            15'd29432: log10_cal = 16'b0000010111010101;
            15'd29433: log10_cal = 16'b0000010111010101;
            15'd29434: log10_cal = 16'b0000010111010101;
            15'd29435: log10_cal = 16'b0000010111010101;
            15'd29436: log10_cal = 16'b0000010111010101;
            15'd29437: log10_cal = 16'b0000010111010101;
            15'd29438: log10_cal = 16'b0000010111010101;
            15'd29439: log10_cal = 16'b0000010111010101;
            15'd29440: log10_cal = 16'b0000010111010101;
            15'd29441: log10_cal = 16'b0000010111010101;
            15'd29442: log10_cal = 16'b0000010111010101;
            15'd29443: log10_cal = 16'b0000010111010101;
            15'd29444: log10_cal = 16'b0000010111010101;
            15'd29445: log10_cal = 16'b0000010111010101;
            15'd29446: log10_cal = 16'b0000010111010101;
            15'd29447: log10_cal = 16'b0000010111010101;
            15'd29448: log10_cal = 16'b0000010111010101;
            15'd29449: log10_cal = 16'b0000010111010101;
            15'd29450: log10_cal = 16'b0000010111010101;
            15'd29451: log10_cal = 16'b0000010111010101;
            15'd29452: log10_cal = 16'b0000010111010101;
            15'd29453: log10_cal = 16'b0000010111010101;
            15'd29454: log10_cal = 16'b0000010111010101;
            15'd29455: log10_cal = 16'b0000010111010101;
            15'd29456: log10_cal = 16'b0000010111010101;
            15'd29457: log10_cal = 16'b0000010111010101;
            15'd29458: log10_cal = 16'b0000010111010101;
            15'd29459: log10_cal = 16'b0000010111010101;
            15'd29460: log10_cal = 16'b0000010111010101;
            15'd29461: log10_cal = 16'b0000010111010101;
            15'd29462: log10_cal = 16'b0000010111010101;
            15'd29463: log10_cal = 16'b0000010111010101;
            15'd29464: log10_cal = 16'b0000010111010110;
            15'd29465: log10_cal = 16'b0000010111010110;
            15'd29466: log10_cal = 16'b0000010111010110;
            15'd29467: log10_cal = 16'b0000010111010110;
            15'd29468: log10_cal = 16'b0000010111010110;
            15'd29469: log10_cal = 16'b0000010111010110;
            15'd29470: log10_cal = 16'b0000010111010110;
            15'd29471: log10_cal = 16'b0000010111010110;
            15'd29472: log10_cal = 16'b0000010111010110;
            15'd29473: log10_cal = 16'b0000010111010110;
            15'd29474: log10_cal = 16'b0000010111010110;
            15'd29475: log10_cal = 16'b0000010111010110;
            15'd29476: log10_cal = 16'b0000010111010110;
            15'd29477: log10_cal = 16'b0000010111010110;
            15'd29478: log10_cal = 16'b0000010111010110;
            15'd29479: log10_cal = 16'b0000010111010110;
            15'd29480: log10_cal = 16'b0000010111010110;
            15'd29481: log10_cal = 16'b0000010111010110;
            15'd29482: log10_cal = 16'b0000010111010110;
            15'd29483: log10_cal = 16'b0000010111010110;
            15'd29484: log10_cal = 16'b0000010111010110;
            15'd29485: log10_cal = 16'b0000010111010110;
            15'd29486: log10_cal = 16'b0000010111010110;
            15'd29487: log10_cal = 16'b0000010111010110;
            15'd29488: log10_cal = 16'b0000010111010110;
            15'd29489: log10_cal = 16'b0000010111010110;
            15'd29490: log10_cal = 16'b0000010111010110;
            15'd29491: log10_cal = 16'b0000010111010110;
            15'd29492: log10_cal = 16'b0000010111010110;
            15'd29493: log10_cal = 16'b0000010111010110;
            15'd29494: log10_cal = 16'b0000010111010110;
            15'd29495: log10_cal = 16'b0000010111010110;
            15'd29496: log10_cal = 16'b0000010111010110;
            15'd29497: log10_cal = 16'b0000010111010110;
            15'd29498: log10_cal = 16'b0000010111010110;
            15'd29499: log10_cal = 16'b0000010111010110;
            15'd29500: log10_cal = 16'b0000010111010110;
            15'd29501: log10_cal = 16'b0000010111010110;
            15'd29502: log10_cal = 16'b0000010111010110;
            15'd29503: log10_cal = 16'b0000010111010110;
            15'd29504: log10_cal = 16'b0000010111010110;
            15'd29505: log10_cal = 16'b0000010111010110;
            15'd29506: log10_cal = 16'b0000010111010110;
            15'd29507: log10_cal = 16'b0000010111010110;
            15'd29508: log10_cal = 16'b0000010111010110;
            15'd29509: log10_cal = 16'b0000010111010110;
            15'd29510: log10_cal = 16'b0000010111010110;
            15'd29511: log10_cal = 16'b0000010111010110;
            15'd29512: log10_cal = 16'b0000010111010110;
            15'd29513: log10_cal = 16'b0000010111010110;
            15'd29514: log10_cal = 16'b0000010111010110;
            15'd29515: log10_cal = 16'b0000010111010110;
            15'd29516: log10_cal = 16'b0000010111010110;
            15'd29517: log10_cal = 16'b0000010111010110;
            15'd29518: log10_cal = 16'b0000010111010110;
            15'd29519: log10_cal = 16'b0000010111010110;
            15'd29520: log10_cal = 16'b0000010111010110;
            15'd29521: log10_cal = 16'b0000010111010110;
            15'd29522: log10_cal = 16'b0000010111010110;
            15'd29523: log10_cal = 16'b0000010111010110;
            15'd29524: log10_cal = 16'b0000010111010110;
            15'd29525: log10_cal = 16'b0000010111010110;
            15'd29526: log10_cal = 16'b0000010111010110;
            15'd29527: log10_cal = 16'b0000010111010110;
            15'd29528: log10_cal = 16'b0000010111010110;
            15'd29529: log10_cal = 16'b0000010111010110;
            15'd29530: log10_cal = 16'b0000010111010111;
            15'd29531: log10_cal = 16'b0000010111010111;
            15'd29532: log10_cal = 16'b0000010111010111;
            15'd29533: log10_cal = 16'b0000010111010111;
            15'd29534: log10_cal = 16'b0000010111010111;
            15'd29535: log10_cal = 16'b0000010111010111;
            15'd29536: log10_cal = 16'b0000010111010111;
            15'd29537: log10_cal = 16'b0000010111010111;
            15'd29538: log10_cal = 16'b0000010111010111;
            15'd29539: log10_cal = 16'b0000010111010111;
            15'd29540: log10_cal = 16'b0000010111010111;
            15'd29541: log10_cal = 16'b0000010111010111;
            15'd29542: log10_cal = 16'b0000010111010111;
            15'd29543: log10_cal = 16'b0000010111010111;
            15'd29544: log10_cal = 16'b0000010111010111;
            15'd29545: log10_cal = 16'b0000010111010111;
            15'd29546: log10_cal = 16'b0000010111010111;
            15'd29547: log10_cal = 16'b0000010111010111;
            15'd29548: log10_cal = 16'b0000010111010111;
            15'd29549: log10_cal = 16'b0000010111010111;
            15'd29550: log10_cal = 16'b0000010111010111;
            15'd29551: log10_cal = 16'b0000010111010111;
            15'd29552: log10_cal = 16'b0000010111010111;
            15'd29553: log10_cal = 16'b0000010111010111;
            15'd29554: log10_cal = 16'b0000010111010111;
            15'd29555: log10_cal = 16'b0000010111010111;
            15'd29556: log10_cal = 16'b0000010111010111;
            15'd29557: log10_cal = 16'b0000010111010111;
            15'd29558: log10_cal = 16'b0000010111010111;
            15'd29559: log10_cal = 16'b0000010111010111;
            15'd29560: log10_cal = 16'b0000010111010111;
            15'd29561: log10_cal = 16'b0000010111010111;
            15'd29562: log10_cal = 16'b0000010111010111;
            15'd29563: log10_cal = 16'b0000010111010111;
            15'd29564: log10_cal = 16'b0000010111010111;
            15'd29565: log10_cal = 16'b0000010111010111;
            15'd29566: log10_cal = 16'b0000010111010111;
            15'd29567: log10_cal = 16'b0000010111010111;
            15'd29568: log10_cal = 16'b0000010111010111;
            15'd29569: log10_cal = 16'b0000010111010111;
            15'd29570: log10_cal = 16'b0000010111010111;
            15'd29571: log10_cal = 16'b0000010111010111;
            15'd29572: log10_cal = 16'b0000010111010111;
            15'd29573: log10_cal = 16'b0000010111010111;
            15'd29574: log10_cal = 16'b0000010111010111;
            15'd29575: log10_cal = 16'b0000010111010111;
            15'd29576: log10_cal = 16'b0000010111010111;
            15'd29577: log10_cal = 16'b0000010111010111;
            15'd29578: log10_cal = 16'b0000010111010111;
            15'd29579: log10_cal = 16'b0000010111010111;
            15'd29580: log10_cal = 16'b0000010111010111;
            15'd29581: log10_cal = 16'b0000010111010111;
            15'd29582: log10_cal = 16'b0000010111010111;
            15'd29583: log10_cal = 16'b0000010111010111;
            15'd29584: log10_cal = 16'b0000010111010111;
            15'd29585: log10_cal = 16'b0000010111010111;
            15'd29586: log10_cal = 16'b0000010111010111;
            15'd29587: log10_cal = 16'b0000010111010111;
            15'd29588: log10_cal = 16'b0000010111010111;
            15'd29589: log10_cal = 16'b0000010111010111;
            15'd29590: log10_cal = 16'b0000010111010111;
            15'd29591: log10_cal = 16'b0000010111010111;
            15'd29592: log10_cal = 16'b0000010111010111;
            15'd29593: log10_cal = 16'b0000010111010111;
            15'd29594: log10_cal = 16'b0000010111010111;
            15'd29595: log10_cal = 16'b0000010111010111;
            15'd29596: log10_cal = 16'b0000010111010111;
            15'd29597: log10_cal = 16'b0000010111011000;
            15'd29598: log10_cal = 16'b0000010111011000;
            15'd29599: log10_cal = 16'b0000010111011000;
            15'd29600: log10_cal = 16'b0000010111011000;
            15'd29601: log10_cal = 16'b0000010111011000;
            15'd29602: log10_cal = 16'b0000010111011000;
            15'd29603: log10_cal = 16'b0000010111011000;
            15'd29604: log10_cal = 16'b0000010111011000;
            15'd29605: log10_cal = 16'b0000010111011000;
            15'd29606: log10_cal = 16'b0000010111011000;
            15'd29607: log10_cal = 16'b0000010111011000;
            15'd29608: log10_cal = 16'b0000010111011000;
            15'd29609: log10_cal = 16'b0000010111011000;
            15'd29610: log10_cal = 16'b0000010111011000;
            15'd29611: log10_cal = 16'b0000010111011000;
            15'd29612: log10_cal = 16'b0000010111011000;
            15'd29613: log10_cal = 16'b0000010111011000;
            15'd29614: log10_cal = 16'b0000010111011000;
            15'd29615: log10_cal = 16'b0000010111011000;
            15'd29616: log10_cal = 16'b0000010111011000;
            15'd29617: log10_cal = 16'b0000010111011000;
            15'd29618: log10_cal = 16'b0000010111011000;
            15'd29619: log10_cal = 16'b0000010111011000;
            15'd29620: log10_cal = 16'b0000010111011000;
            15'd29621: log10_cal = 16'b0000010111011000;
            15'd29622: log10_cal = 16'b0000010111011000;
            15'd29623: log10_cal = 16'b0000010111011000;
            15'd29624: log10_cal = 16'b0000010111011000;
            15'd29625: log10_cal = 16'b0000010111011000;
            15'd29626: log10_cal = 16'b0000010111011000;
            15'd29627: log10_cal = 16'b0000010111011000;
            15'd29628: log10_cal = 16'b0000010111011000;
            15'd29629: log10_cal = 16'b0000010111011000;
            15'd29630: log10_cal = 16'b0000010111011000;
            15'd29631: log10_cal = 16'b0000010111011000;
            15'd29632: log10_cal = 16'b0000010111011000;
            15'd29633: log10_cal = 16'b0000010111011000;
            15'd29634: log10_cal = 16'b0000010111011000;
            15'd29635: log10_cal = 16'b0000010111011000;
            15'd29636: log10_cal = 16'b0000010111011000;
            15'd29637: log10_cal = 16'b0000010111011000;
            15'd29638: log10_cal = 16'b0000010111011000;
            15'd29639: log10_cal = 16'b0000010111011000;
            15'd29640: log10_cal = 16'b0000010111011000;
            15'd29641: log10_cal = 16'b0000010111011000;
            15'd29642: log10_cal = 16'b0000010111011000;
            15'd29643: log10_cal = 16'b0000010111011000;
            15'd29644: log10_cal = 16'b0000010111011000;
            15'd29645: log10_cal = 16'b0000010111011000;
            15'd29646: log10_cal = 16'b0000010111011000;
            15'd29647: log10_cal = 16'b0000010111011000;
            15'd29648: log10_cal = 16'b0000010111011000;
            15'd29649: log10_cal = 16'b0000010111011000;
            15'd29650: log10_cal = 16'b0000010111011000;
            15'd29651: log10_cal = 16'b0000010111011000;
            15'd29652: log10_cal = 16'b0000010111011000;
            15'd29653: log10_cal = 16'b0000010111011000;
            15'd29654: log10_cal = 16'b0000010111011000;
            15'd29655: log10_cal = 16'b0000010111011000;
            15'd29656: log10_cal = 16'b0000010111011000;
            15'd29657: log10_cal = 16'b0000010111011000;
            15'd29658: log10_cal = 16'b0000010111011000;
            15'd29659: log10_cal = 16'b0000010111011000;
            15'd29660: log10_cal = 16'b0000010111011000;
            15'd29661: log10_cal = 16'b0000010111011000;
            15'd29662: log10_cal = 16'b0000010111011000;
            15'd29663: log10_cal = 16'b0000010111011001;
            15'd29664: log10_cal = 16'b0000010111011001;
            15'd29665: log10_cal = 16'b0000010111011001;
            15'd29666: log10_cal = 16'b0000010111011001;
            15'd29667: log10_cal = 16'b0000010111011001;
            15'd29668: log10_cal = 16'b0000010111011001;
            15'd29669: log10_cal = 16'b0000010111011001;
            15'd29670: log10_cal = 16'b0000010111011001;
            15'd29671: log10_cal = 16'b0000010111011001;
            15'd29672: log10_cal = 16'b0000010111011001;
            15'd29673: log10_cal = 16'b0000010111011001;
            15'd29674: log10_cal = 16'b0000010111011001;
            15'd29675: log10_cal = 16'b0000010111011001;
            15'd29676: log10_cal = 16'b0000010111011001;
            15'd29677: log10_cal = 16'b0000010111011001;
            15'd29678: log10_cal = 16'b0000010111011001;
            15'd29679: log10_cal = 16'b0000010111011001;
            15'd29680: log10_cal = 16'b0000010111011001;
            15'd29681: log10_cal = 16'b0000010111011001;
            15'd29682: log10_cal = 16'b0000010111011001;
            15'd29683: log10_cal = 16'b0000010111011001;
            15'd29684: log10_cal = 16'b0000010111011001;
            15'd29685: log10_cal = 16'b0000010111011001;
            15'd29686: log10_cal = 16'b0000010111011001;
            15'd29687: log10_cal = 16'b0000010111011001;
            15'd29688: log10_cal = 16'b0000010111011001;
            15'd29689: log10_cal = 16'b0000010111011001;
            15'd29690: log10_cal = 16'b0000010111011001;
            15'd29691: log10_cal = 16'b0000010111011001;
            15'd29692: log10_cal = 16'b0000010111011001;
            15'd29693: log10_cal = 16'b0000010111011001;
            15'd29694: log10_cal = 16'b0000010111011001;
            15'd29695: log10_cal = 16'b0000010111011001;
            15'd29696: log10_cal = 16'b0000010111011001;
            15'd29697: log10_cal = 16'b0000010111011001;
            15'd29698: log10_cal = 16'b0000010111011001;
            15'd29699: log10_cal = 16'b0000010111011001;
            15'd29700: log10_cal = 16'b0000010111011001;
            15'd29701: log10_cal = 16'b0000010111011001;
            15'd29702: log10_cal = 16'b0000010111011001;
            15'd29703: log10_cal = 16'b0000010111011001;
            15'd29704: log10_cal = 16'b0000010111011001;
            15'd29705: log10_cal = 16'b0000010111011001;
            15'd29706: log10_cal = 16'b0000010111011001;
            15'd29707: log10_cal = 16'b0000010111011001;
            15'd29708: log10_cal = 16'b0000010111011001;
            15'd29709: log10_cal = 16'b0000010111011001;
            15'd29710: log10_cal = 16'b0000010111011001;
            15'd29711: log10_cal = 16'b0000010111011001;
            15'd29712: log10_cal = 16'b0000010111011001;
            15'd29713: log10_cal = 16'b0000010111011001;
            15'd29714: log10_cal = 16'b0000010111011001;
            15'd29715: log10_cal = 16'b0000010111011001;
            15'd29716: log10_cal = 16'b0000010111011001;
            15'd29717: log10_cal = 16'b0000010111011001;
            15'd29718: log10_cal = 16'b0000010111011001;
            15'd29719: log10_cal = 16'b0000010111011001;
            15'd29720: log10_cal = 16'b0000010111011001;
            15'd29721: log10_cal = 16'b0000010111011001;
            15'd29722: log10_cal = 16'b0000010111011001;
            15'd29723: log10_cal = 16'b0000010111011001;
            15'd29724: log10_cal = 16'b0000010111011001;
            15'd29725: log10_cal = 16'b0000010111011001;
            15'd29726: log10_cal = 16'b0000010111011001;
            15'd29727: log10_cal = 16'b0000010111011001;
            15'd29728: log10_cal = 16'b0000010111011001;
            15'd29729: log10_cal = 16'b0000010111011001;
            15'd29730: log10_cal = 16'b0000010111011010;
            15'd29731: log10_cal = 16'b0000010111011010;
            15'd29732: log10_cal = 16'b0000010111011010;
            15'd29733: log10_cal = 16'b0000010111011010;
            15'd29734: log10_cal = 16'b0000010111011010;
            15'd29735: log10_cal = 16'b0000010111011010;
            15'd29736: log10_cal = 16'b0000010111011010;
            15'd29737: log10_cal = 16'b0000010111011010;
            15'd29738: log10_cal = 16'b0000010111011010;
            15'd29739: log10_cal = 16'b0000010111011010;
            15'd29740: log10_cal = 16'b0000010111011010;
            15'd29741: log10_cal = 16'b0000010111011010;
            15'd29742: log10_cal = 16'b0000010111011010;
            15'd29743: log10_cal = 16'b0000010111011010;
            15'd29744: log10_cal = 16'b0000010111011010;
            15'd29745: log10_cal = 16'b0000010111011010;
            15'd29746: log10_cal = 16'b0000010111011010;
            15'd29747: log10_cal = 16'b0000010111011010;
            15'd29748: log10_cal = 16'b0000010111011010;
            15'd29749: log10_cal = 16'b0000010111011010;
            15'd29750: log10_cal = 16'b0000010111011010;
            15'd29751: log10_cal = 16'b0000010111011010;
            15'd29752: log10_cal = 16'b0000010111011010;
            15'd29753: log10_cal = 16'b0000010111011010;
            15'd29754: log10_cal = 16'b0000010111011010;
            15'd29755: log10_cal = 16'b0000010111011010;
            15'd29756: log10_cal = 16'b0000010111011010;
            15'd29757: log10_cal = 16'b0000010111011010;
            15'd29758: log10_cal = 16'b0000010111011010;
            15'd29759: log10_cal = 16'b0000010111011010;
            15'd29760: log10_cal = 16'b0000010111011010;
            15'd29761: log10_cal = 16'b0000010111011010;
            15'd29762: log10_cal = 16'b0000010111011010;
            15'd29763: log10_cal = 16'b0000010111011010;
            15'd29764: log10_cal = 16'b0000010111011010;
            15'd29765: log10_cal = 16'b0000010111011010;
            15'd29766: log10_cal = 16'b0000010111011010;
            15'd29767: log10_cal = 16'b0000010111011010;
            15'd29768: log10_cal = 16'b0000010111011010;
            15'd29769: log10_cal = 16'b0000010111011010;
            15'd29770: log10_cal = 16'b0000010111011010;
            15'd29771: log10_cal = 16'b0000010111011010;
            15'd29772: log10_cal = 16'b0000010111011010;
            15'd29773: log10_cal = 16'b0000010111011010;
            15'd29774: log10_cal = 16'b0000010111011010;
            15'd29775: log10_cal = 16'b0000010111011010;
            15'd29776: log10_cal = 16'b0000010111011010;
            15'd29777: log10_cal = 16'b0000010111011010;
            15'd29778: log10_cal = 16'b0000010111011010;
            15'd29779: log10_cal = 16'b0000010111011010;
            15'd29780: log10_cal = 16'b0000010111011010;
            15'd29781: log10_cal = 16'b0000010111011010;
            15'd29782: log10_cal = 16'b0000010111011010;
            15'd29783: log10_cal = 16'b0000010111011010;
            15'd29784: log10_cal = 16'b0000010111011010;
            15'd29785: log10_cal = 16'b0000010111011010;
            15'd29786: log10_cal = 16'b0000010111011010;
            15'd29787: log10_cal = 16'b0000010111011010;
            15'd29788: log10_cal = 16'b0000010111011010;
            15'd29789: log10_cal = 16'b0000010111011010;
            15'd29790: log10_cal = 16'b0000010111011010;
            15'd29791: log10_cal = 16'b0000010111011010;
            15'd29792: log10_cal = 16'b0000010111011010;
            15'd29793: log10_cal = 16'b0000010111011010;
            15'd29794: log10_cal = 16'b0000010111011010;
            15'd29795: log10_cal = 16'b0000010111011010;
            15'd29796: log10_cal = 16'b0000010111011010;
            15'd29797: log10_cal = 16'b0000010111011011;
            15'd29798: log10_cal = 16'b0000010111011011;
            15'd29799: log10_cal = 16'b0000010111011011;
            15'd29800: log10_cal = 16'b0000010111011011;
            15'd29801: log10_cal = 16'b0000010111011011;
            15'd29802: log10_cal = 16'b0000010111011011;
            15'd29803: log10_cal = 16'b0000010111011011;
            15'd29804: log10_cal = 16'b0000010111011011;
            15'd29805: log10_cal = 16'b0000010111011011;
            15'd29806: log10_cal = 16'b0000010111011011;
            15'd29807: log10_cal = 16'b0000010111011011;
            15'd29808: log10_cal = 16'b0000010111011011;
            15'd29809: log10_cal = 16'b0000010111011011;
            15'd29810: log10_cal = 16'b0000010111011011;
            15'd29811: log10_cal = 16'b0000010111011011;
            15'd29812: log10_cal = 16'b0000010111011011;
            15'd29813: log10_cal = 16'b0000010111011011;
            15'd29814: log10_cal = 16'b0000010111011011;
            15'd29815: log10_cal = 16'b0000010111011011;
            15'd29816: log10_cal = 16'b0000010111011011;
            15'd29817: log10_cal = 16'b0000010111011011;
            15'd29818: log10_cal = 16'b0000010111011011;
            15'd29819: log10_cal = 16'b0000010111011011;
            15'd29820: log10_cal = 16'b0000010111011011;
            15'd29821: log10_cal = 16'b0000010111011011;
            15'd29822: log10_cal = 16'b0000010111011011;
            15'd29823: log10_cal = 16'b0000010111011011;
            15'd29824: log10_cal = 16'b0000010111011011;
            15'd29825: log10_cal = 16'b0000010111011011;
            15'd29826: log10_cal = 16'b0000010111011011;
            15'd29827: log10_cal = 16'b0000010111011011;
            15'd29828: log10_cal = 16'b0000010111011011;
            15'd29829: log10_cal = 16'b0000010111011011;
            15'd29830: log10_cal = 16'b0000010111011011;
            15'd29831: log10_cal = 16'b0000010111011011;
            15'd29832: log10_cal = 16'b0000010111011011;
            15'd29833: log10_cal = 16'b0000010111011011;
            15'd29834: log10_cal = 16'b0000010111011011;
            15'd29835: log10_cal = 16'b0000010111011011;
            15'd29836: log10_cal = 16'b0000010111011011;
            15'd29837: log10_cal = 16'b0000010111011011;
            15'd29838: log10_cal = 16'b0000010111011011;
            15'd29839: log10_cal = 16'b0000010111011011;
            15'd29840: log10_cal = 16'b0000010111011011;
            15'd29841: log10_cal = 16'b0000010111011011;
            15'd29842: log10_cal = 16'b0000010111011011;
            15'd29843: log10_cal = 16'b0000010111011011;
            15'd29844: log10_cal = 16'b0000010111011011;
            15'd29845: log10_cal = 16'b0000010111011011;
            15'd29846: log10_cal = 16'b0000010111011011;
            15'd29847: log10_cal = 16'b0000010111011011;
            15'd29848: log10_cal = 16'b0000010111011011;
            15'd29849: log10_cal = 16'b0000010111011011;
            15'd29850: log10_cal = 16'b0000010111011011;
            15'd29851: log10_cal = 16'b0000010111011011;
            15'd29852: log10_cal = 16'b0000010111011011;
            15'd29853: log10_cal = 16'b0000010111011011;
            15'd29854: log10_cal = 16'b0000010111011011;
            15'd29855: log10_cal = 16'b0000010111011011;
            15'd29856: log10_cal = 16'b0000010111011011;
            15'd29857: log10_cal = 16'b0000010111011011;
            15'd29858: log10_cal = 16'b0000010111011011;
            15'd29859: log10_cal = 16'b0000010111011011;
            15'd29860: log10_cal = 16'b0000010111011011;
            15'd29861: log10_cal = 16'b0000010111011011;
            15'd29862: log10_cal = 16'b0000010111011011;
            15'd29863: log10_cal = 16'b0000010111011011;
            15'd29864: log10_cal = 16'b0000010111011100;
            15'd29865: log10_cal = 16'b0000010111011100;
            15'd29866: log10_cal = 16'b0000010111011100;
            15'd29867: log10_cal = 16'b0000010111011100;
            15'd29868: log10_cal = 16'b0000010111011100;
            15'd29869: log10_cal = 16'b0000010111011100;
            15'd29870: log10_cal = 16'b0000010111011100;
            15'd29871: log10_cal = 16'b0000010111011100;
            15'd29872: log10_cal = 16'b0000010111011100;
            15'd29873: log10_cal = 16'b0000010111011100;
            15'd29874: log10_cal = 16'b0000010111011100;
            15'd29875: log10_cal = 16'b0000010111011100;
            15'd29876: log10_cal = 16'b0000010111011100;
            15'd29877: log10_cal = 16'b0000010111011100;
            15'd29878: log10_cal = 16'b0000010111011100;
            15'd29879: log10_cal = 16'b0000010111011100;
            15'd29880: log10_cal = 16'b0000010111011100;
            15'd29881: log10_cal = 16'b0000010111011100;
            15'd29882: log10_cal = 16'b0000010111011100;
            15'd29883: log10_cal = 16'b0000010111011100;
            15'd29884: log10_cal = 16'b0000010111011100;
            15'd29885: log10_cal = 16'b0000010111011100;
            15'd29886: log10_cal = 16'b0000010111011100;
            15'd29887: log10_cal = 16'b0000010111011100;
            15'd29888: log10_cal = 16'b0000010111011100;
            15'd29889: log10_cal = 16'b0000010111011100;
            15'd29890: log10_cal = 16'b0000010111011100;
            15'd29891: log10_cal = 16'b0000010111011100;
            15'd29892: log10_cal = 16'b0000010111011100;
            15'd29893: log10_cal = 16'b0000010111011100;
            15'd29894: log10_cal = 16'b0000010111011100;
            15'd29895: log10_cal = 16'b0000010111011100;
            15'd29896: log10_cal = 16'b0000010111011100;
            15'd29897: log10_cal = 16'b0000010111011100;
            15'd29898: log10_cal = 16'b0000010111011100;
            15'd29899: log10_cal = 16'b0000010111011100;
            15'd29900: log10_cal = 16'b0000010111011100;
            15'd29901: log10_cal = 16'b0000010111011100;
            15'd29902: log10_cal = 16'b0000010111011100;
            15'd29903: log10_cal = 16'b0000010111011100;
            15'd29904: log10_cal = 16'b0000010111011100;
            15'd29905: log10_cal = 16'b0000010111011100;
            15'd29906: log10_cal = 16'b0000010111011100;
            15'd29907: log10_cal = 16'b0000010111011100;
            15'd29908: log10_cal = 16'b0000010111011100;
            15'd29909: log10_cal = 16'b0000010111011100;
            15'd29910: log10_cal = 16'b0000010111011100;
            15'd29911: log10_cal = 16'b0000010111011100;
            15'd29912: log10_cal = 16'b0000010111011100;
            15'd29913: log10_cal = 16'b0000010111011100;
            15'd29914: log10_cal = 16'b0000010111011100;
            15'd29915: log10_cal = 16'b0000010111011100;
            15'd29916: log10_cal = 16'b0000010111011100;
            15'd29917: log10_cal = 16'b0000010111011100;
            15'd29918: log10_cal = 16'b0000010111011100;
            15'd29919: log10_cal = 16'b0000010111011100;
            15'd29920: log10_cal = 16'b0000010111011100;
            15'd29921: log10_cal = 16'b0000010111011100;
            15'd29922: log10_cal = 16'b0000010111011100;
            15'd29923: log10_cal = 16'b0000010111011100;
            15'd29924: log10_cal = 16'b0000010111011100;
            15'd29925: log10_cal = 16'b0000010111011100;
            15'd29926: log10_cal = 16'b0000010111011100;
            15'd29927: log10_cal = 16'b0000010111011100;
            15'd29928: log10_cal = 16'b0000010111011100;
            15'd29929: log10_cal = 16'b0000010111011100;
            15'd29930: log10_cal = 16'b0000010111011100;
            15'd29931: log10_cal = 16'b0000010111011101;
            15'd29932: log10_cal = 16'b0000010111011101;
            15'd29933: log10_cal = 16'b0000010111011101;
            15'd29934: log10_cal = 16'b0000010111011101;
            15'd29935: log10_cal = 16'b0000010111011101;
            15'd29936: log10_cal = 16'b0000010111011101;
            15'd29937: log10_cal = 16'b0000010111011101;
            15'd29938: log10_cal = 16'b0000010111011101;
            15'd29939: log10_cal = 16'b0000010111011101;
            15'd29940: log10_cal = 16'b0000010111011101;
            15'd29941: log10_cal = 16'b0000010111011101;
            15'd29942: log10_cal = 16'b0000010111011101;
            15'd29943: log10_cal = 16'b0000010111011101;
            15'd29944: log10_cal = 16'b0000010111011101;
            15'd29945: log10_cal = 16'b0000010111011101;
            15'd29946: log10_cal = 16'b0000010111011101;
            15'd29947: log10_cal = 16'b0000010111011101;
            15'd29948: log10_cal = 16'b0000010111011101;
            15'd29949: log10_cal = 16'b0000010111011101;
            15'd29950: log10_cal = 16'b0000010111011101;
            15'd29951: log10_cal = 16'b0000010111011101;
            15'd29952: log10_cal = 16'b0000010111011101;
            15'd29953: log10_cal = 16'b0000010111011101;
            15'd29954: log10_cal = 16'b0000010111011101;
            15'd29955: log10_cal = 16'b0000010111011101;
            15'd29956: log10_cal = 16'b0000010111011101;
            15'd29957: log10_cal = 16'b0000010111011101;
            15'd29958: log10_cal = 16'b0000010111011101;
            15'd29959: log10_cal = 16'b0000010111011101;
            15'd29960: log10_cal = 16'b0000010111011101;
            15'd29961: log10_cal = 16'b0000010111011101;
            15'd29962: log10_cal = 16'b0000010111011101;
            15'd29963: log10_cal = 16'b0000010111011101;
            15'd29964: log10_cal = 16'b0000010111011101;
            15'd29965: log10_cal = 16'b0000010111011101;
            15'd29966: log10_cal = 16'b0000010111011101;
            15'd29967: log10_cal = 16'b0000010111011101;
            15'd29968: log10_cal = 16'b0000010111011101;
            15'd29969: log10_cal = 16'b0000010111011101;
            15'd29970: log10_cal = 16'b0000010111011101;
            15'd29971: log10_cal = 16'b0000010111011101;
            15'd29972: log10_cal = 16'b0000010111011101;
            15'd29973: log10_cal = 16'b0000010111011101;
            15'd29974: log10_cal = 16'b0000010111011101;
            15'd29975: log10_cal = 16'b0000010111011101;
            15'd29976: log10_cal = 16'b0000010111011101;
            15'd29977: log10_cal = 16'b0000010111011101;
            15'd29978: log10_cal = 16'b0000010111011101;
            15'd29979: log10_cal = 16'b0000010111011101;
            15'd29980: log10_cal = 16'b0000010111011101;
            15'd29981: log10_cal = 16'b0000010111011101;
            15'd29982: log10_cal = 16'b0000010111011101;
            15'd29983: log10_cal = 16'b0000010111011101;
            15'd29984: log10_cal = 16'b0000010111011101;
            15'd29985: log10_cal = 16'b0000010111011101;
            15'd29986: log10_cal = 16'b0000010111011101;
            15'd29987: log10_cal = 16'b0000010111011101;
            15'd29988: log10_cal = 16'b0000010111011101;
            15'd29989: log10_cal = 16'b0000010111011101;
            15'd29990: log10_cal = 16'b0000010111011101;
            15'd29991: log10_cal = 16'b0000010111011101;
            15'd29992: log10_cal = 16'b0000010111011101;
            15'd29993: log10_cal = 16'b0000010111011101;
            15'd29994: log10_cal = 16'b0000010111011101;
            15'd29995: log10_cal = 16'b0000010111011101;
            15'd29996: log10_cal = 16'b0000010111011101;
            15'd29997: log10_cal = 16'b0000010111011101;
            15'd29998: log10_cal = 16'b0000010111011101;
            15'd29999: log10_cal = 16'b0000010111011110;
            15'd30000: log10_cal = 16'b0000010111011110;
            15'd30001: log10_cal = 16'b0000010111011110;
            15'd30002: log10_cal = 16'b0000010111011110;
            15'd30003: log10_cal = 16'b0000010111011110;
            15'd30004: log10_cal = 16'b0000010111011110;
            15'd30005: log10_cal = 16'b0000010111011110;
            15'd30006: log10_cal = 16'b0000010111011110;
            15'd30007: log10_cal = 16'b0000010111011110;
            15'd30008: log10_cal = 16'b0000010111011110;
            15'd30009: log10_cal = 16'b0000010111011110;
            15'd30010: log10_cal = 16'b0000010111011110;
            15'd30011: log10_cal = 16'b0000010111011110;
            15'd30012: log10_cal = 16'b0000010111011110;
            15'd30013: log10_cal = 16'b0000010111011110;
            15'd30014: log10_cal = 16'b0000010111011110;
            15'd30015: log10_cal = 16'b0000010111011110;
            15'd30016: log10_cal = 16'b0000010111011110;
            15'd30017: log10_cal = 16'b0000010111011110;
            15'd30018: log10_cal = 16'b0000010111011110;
            15'd30019: log10_cal = 16'b0000010111011110;
            15'd30020: log10_cal = 16'b0000010111011110;
            15'd30021: log10_cal = 16'b0000010111011110;
            15'd30022: log10_cal = 16'b0000010111011110;
            15'd30023: log10_cal = 16'b0000010111011110;
            15'd30024: log10_cal = 16'b0000010111011110;
            15'd30025: log10_cal = 16'b0000010111011110;
            15'd30026: log10_cal = 16'b0000010111011110;
            15'd30027: log10_cal = 16'b0000010111011110;
            15'd30028: log10_cal = 16'b0000010111011110;
            15'd30029: log10_cal = 16'b0000010111011110;
            15'd30030: log10_cal = 16'b0000010111011110;
            15'd30031: log10_cal = 16'b0000010111011110;
            15'd30032: log10_cal = 16'b0000010111011110;
            15'd30033: log10_cal = 16'b0000010111011110;
            15'd30034: log10_cal = 16'b0000010111011110;
            15'd30035: log10_cal = 16'b0000010111011110;
            15'd30036: log10_cal = 16'b0000010111011110;
            15'd30037: log10_cal = 16'b0000010111011110;
            15'd30038: log10_cal = 16'b0000010111011110;
            15'd30039: log10_cal = 16'b0000010111011110;
            15'd30040: log10_cal = 16'b0000010111011110;
            15'd30041: log10_cal = 16'b0000010111011110;
            15'd30042: log10_cal = 16'b0000010111011110;
            15'd30043: log10_cal = 16'b0000010111011110;
            15'd30044: log10_cal = 16'b0000010111011110;
            15'd30045: log10_cal = 16'b0000010111011110;
            15'd30046: log10_cal = 16'b0000010111011110;
            15'd30047: log10_cal = 16'b0000010111011110;
            15'd30048: log10_cal = 16'b0000010111011110;
            15'd30049: log10_cal = 16'b0000010111011110;
            15'd30050: log10_cal = 16'b0000010111011110;
            15'd30051: log10_cal = 16'b0000010111011110;
            15'd30052: log10_cal = 16'b0000010111011110;
            15'd30053: log10_cal = 16'b0000010111011110;
            15'd30054: log10_cal = 16'b0000010111011110;
            15'd30055: log10_cal = 16'b0000010111011110;
            15'd30056: log10_cal = 16'b0000010111011110;
            15'd30057: log10_cal = 16'b0000010111011110;
            15'd30058: log10_cal = 16'b0000010111011110;
            15'd30059: log10_cal = 16'b0000010111011110;
            15'd30060: log10_cal = 16'b0000010111011110;
            15'd30061: log10_cal = 16'b0000010111011110;
            15'd30062: log10_cal = 16'b0000010111011110;
            15'd30063: log10_cal = 16'b0000010111011110;
            15'd30064: log10_cal = 16'b0000010111011110;
            15'd30065: log10_cal = 16'b0000010111011110;
            15'd30066: log10_cal = 16'b0000010111011111;
            15'd30067: log10_cal = 16'b0000010111011111;
            15'd30068: log10_cal = 16'b0000010111011111;
            15'd30069: log10_cal = 16'b0000010111011111;
            15'd30070: log10_cal = 16'b0000010111011111;
            15'd30071: log10_cal = 16'b0000010111011111;
            15'd30072: log10_cal = 16'b0000010111011111;
            15'd30073: log10_cal = 16'b0000010111011111;
            15'd30074: log10_cal = 16'b0000010111011111;
            15'd30075: log10_cal = 16'b0000010111011111;
            15'd30076: log10_cal = 16'b0000010111011111;
            15'd30077: log10_cal = 16'b0000010111011111;
            15'd30078: log10_cal = 16'b0000010111011111;
            15'd30079: log10_cal = 16'b0000010111011111;
            15'd30080: log10_cal = 16'b0000010111011111;
            15'd30081: log10_cal = 16'b0000010111011111;
            15'd30082: log10_cal = 16'b0000010111011111;
            15'd30083: log10_cal = 16'b0000010111011111;
            15'd30084: log10_cal = 16'b0000010111011111;
            15'd30085: log10_cal = 16'b0000010111011111;
            15'd30086: log10_cal = 16'b0000010111011111;
            15'd30087: log10_cal = 16'b0000010111011111;
            15'd30088: log10_cal = 16'b0000010111011111;
            15'd30089: log10_cal = 16'b0000010111011111;
            15'd30090: log10_cal = 16'b0000010111011111;
            15'd30091: log10_cal = 16'b0000010111011111;
            15'd30092: log10_cal = 16'b0000010111011111;
            15'd30093: log10_cal = 16'b0000010111011111;
            15'd30094: log10_cal = 16'b0000010111011111;
            15'd30095: log10_cal = 16'b0000010111011111;
            15'd30096: log10_cal = 16'b0000010111011111;
            15'd30097: log10_cal = 16'b0000010111011111;
            15'd30098: log10_cal = 16'b0000010111011111;
            15'd30099: log10_cal = 16'b0000010111011111;
            15'd30100: log10_cal = 16'b0000010111011111;
            15'd30101: log10_cal = 16'b0000010111011111;
            15'd30102: log10_cal = 16'b0000010111011111;
            15'd30103: log10_cal = 16'b0000010111011111;
            15'd30104: log10_cal = 16'b0000010111011111;
            15'd30105: log10_cal = 16'b0000010111011111;
            15'd30106: log10_cal = 16'b0000010111011111;
            15'd30107: log10_cal = 16'b0000010111011111;
            15'd30108: log10_cal = 16'b0000010111011111;
            15'd30109: log10_cal = 16'b0000010111011111;
            15'd30110: log10_cal = 16'b0000010111011111;
            15'd30111: log10_cal = 16'b0000010111011111;
            15'd30112: log10_cal = 16'b0000010111011111;
            15'd30113: log10_cal = 16'b0000010111011111;
            15'd30114: log10_cal = 16'b0000010111011111;
            15'd30115: log10_cal = 16'b0000010111011111;
            15'd30116: log10_cal = 16'b0000010111011111;
            15'd30117: log10_cal = 16'b0000010111011111;
            15'd30118: log10_cal = 16'b0000010111011111;
            15'd30119: log10_cal = 16'b0000010111011111;
            15'd30120: log10_cal = 16'b0000010111011111;
            15'd30121: log10_cal = 16'b0000010111011111;
            15'd30122: log10_cal = 16'b0000010111011111;
            15'd30123: log10_cal = 16'b0000010111011111;
            15'd30124: log10_cal = 16'b0000010111011111;
            15'd30125: log10_cal = 16'b0000010111011111;
            15'd30126: log10_cal = 16'b0000010111011111;
            15'd30127: log10_cal = 16'b0000010111011111;
            15'd30128: log10_cal = 16'b0000010111011111;
            15'd30129: log10_cal = 16'b0000010111011111;
            15'd30130: log10_cal = 16'b0000010111011111;
            15'd30131: log10_cal = 16'b0000010111011111;
            15'd30132: log10_cal = 16'b0000010111011111;
            15'd30133: log10_cal = 16'b0000010111011111;
            15'd30134: log10_cal = 16'b0000010111100000;
            15'd30135: log10_cal = 16'b0000010111100000;
            15'd30136: log10_cal = 16'b0000010111100000;
            15'd30137: log10_cal = 16'b0000010111100000;
            15'd30138: log10_cal = 16'b0000010111100000;
            15'd30139: log10_cal = 16'b0000010111100000;
            15'd30140: log10_cal = 16'b0000010111100000;
            15'd30141: log10_cal = 16'b0000010111100000;
            15'd30142: log10_cal = 16'b0000010111100000;
            15'd30143: log10_cal = 16'b0000010111100000;
            15'd30144: log10_cal = 16'b0000010111100000;
            15'd30145: log10_cal = 16'b0000010111100000;
            15'd30146: log10_cal = 16'b0000010111100000;
            15'd30147: log10_cal = 16'b0000010111100000;
            15'd30148: log10_cal = 16'b0000010111100000;
            15'd30149: log10_cal = 16'b0000010111100000;
            15'd30150: log10_cal = 16'b0000010111100000;
            15'd30151: log10_cal = 16'b0000010111100000;
            15'd30152: log10_cal = 16'b0000010111100000;
            15'd30153: log10_cal = 16'b0000010111100000;
            15'd30154: log10_cal = 16'b0000010111100000;
            15'd30155: log10_cal = 16'b0000010111100000;
            15'd30156: log10_cal = 16'b0000010111100000;
            15'd30157: log10_cal = 16'b0000010111100000;
            15'd30158: log10_cal = 16'b0000010111100000;
            15'd30159: log10_cal = 16'b0000010111100000;
            15'd30160: log10_cal = 16'b0000010111100000;
            15'd30161: log10_cal = 16'b0000010111100000;
            15'd30162: log10_cal = 16'b0000010111100000;
            15'd30163: log10_cal = 16'b0000010111100000;
            15'd30164: log10_cal = 16'b0000010111100000;
            15'd30165: log10_cal = 16'b0000010111100000;
            15'd30166: log10_cal = 16'b0000010111100000;
            15'd30167: log10_cal = 16'b0000010111100000;
            15'd30168: log10_cal = 16'b0000010111100000;
            15'd30169: log10_cal = 16'b0000010111100000;
            15'd30170: log10_cal = 16'b0000010111100000;
            15'd30171: log10_cal = 16'b0000010111100000;
            15'd30172: log10_cal = 16'b0000010111100000;
            15'd30173: log10_cal = 16'b0000010111100000;
            15'd30174: log10_cal = 16'b0000010111100000;
            15'd30175: log10_cal = 16'b0000010111100000;
            15'd30176: log10_cal = 16'b0000010111100000;
            15'd30177: log10_cal = 16'b0000010111100000;
            15'd30178: log10_cal = 16'b0000010111100000;
            15'd30179: log10_cal = 16'b0000010111100000;
            15'd30180: log10_cal = 16'b0000010111100000;
            15'd30181: log10_cal = 16'b0000010111100000;
            15'd30182: log10_cal = 16'b0000010111100000;
            15'd30183: log10_cal = 16'b0000010111100000;
            15'd30184: log10_cal = 16'b0000010111100000;
            15'd30185: log10_cal = 16'b0000010111100000;
            15'd30186: log10_cal = 16'b0000010111100000;
            15'd30187: log10_cal = 16'b0000010111100000;
            15'd30188: log10_cal = 16'b0000010111100000;
            15'd30189: log10_cal = 16'b0000010111100000;
            15'd30190: log10_cal = 16'b0000010111100000;
            15'd30191: log10_cal = 16'b0000010111100000;
            15'd30192: log10_cal = 16'b0000010111100000;
            15'd30193: log10_cal = 16'b0000010111100000;
            15'd30194: log10_cal = 16'b0000010111100000;
            15'd30195: log10_cal = 16'b0000010111100000;
            15'd30196: log10_cal = 16'b0000010111100000;
            15'd30197: log10_cal = 16'b0000010111100000;
            15'd30198: log10_cal = 16'b0000010111100000;
            15'd30199: log10_cal = 16'b0000010111100000;
            15'd30200: log10_cal = 16'b0000010111100000;
            15'd30201: log10_cal = 16'b0000010111100000;
            15'd30202: log10_cal = 16'b0000010111100001;
            15'd30203: log10_cal = 16'b0000010111100001;
            15'd30204: log10_cal = 16'b0000010111100001;
            15'd30205: log10_cal = 16'b0000010111100001;
            15'd30206: log10_cal = 16'b0000010111100001;
            15'd30207: log10_cal = 16'b0000010111100001;
            15'd30208: log10_cal = 16'b0000010111100001;
            15'd30209: log10_cal = 16'b0000010111100001;
            15'd30210: log10_cal = 16'b0000010111100001;
            15'd30211: log10_cal = 16'b0000010111100001;
            15'd30212: log10_cal = 16'b0000010111100001;
            15'd30213: log10_cal = 16'b0000010111100001;
            15'd30214: log10_cal = 16'b0000010111100001;
            15'd30215: log10_cal = 16'b0000010111100001;
            15'd30216: log10_cal = 16'b0000010111100001;
            15'd30217: log10_cal = 16'b0000010111100001;
            15'd30218: log10_cal = 16'b0000010111100001;
            15'd30219: log10_cal = 16'b0000010111100001;
            15'd30220: log10_cal = 16'b0000010111100001;
            15'd30221: log10_cal = 16'b0000010111100001;
            15'd30222: log10_cal = 16'b0000010111100001;
            15'd30223: log10_cal = 16'b0000010111100001;
            15'd30224: log10_cal = 16'b0000010111100001;
            15'd30225: log10_cal = 16'b0000010111100001;
            15'd30226: log10_cal = 16'b0000010111100001;
            15'd30227: log10_cal = 16'b0000010111100001;
            15'd30228: log10_cal = 16'b0000010111100001;
            15'd30229: log10_cal = 16'b0000010111100001;
            15'd30230: log10_cal = 16'b0000010111100001;
            15'd30231: log10_cal = 16'b0000010111100001;
            15'd30232: log10_cal = 16'b0000010111100001;
            15'd30233: log10_cal = 16'b0000010111100001;
            15'd30234: log10_cal = 16'b0000010111100001;
            15'd30235: log10_cal = 16'b0000010111100001;
            15'd30236: log10_cal = 16'b0000010111100001;
            15'd30237: log10_cal = 16'b0000010111100001;
            15'd30238: log10_cal = 16'b0000010111100001;
            15'd30239: log10_cal = 16'b0000010111100001;
            15'd30240: log10_cal = 16'b0000010111100001;
            15'd30241: log10_cal = 16'b0000010111100001;
            15'd30242: log10_cal = 16'b0000010111100001;
            15'd30243: log10_cal = 16'b0000010111100001;
            15'd30244: log10_cal = 16'b0000010111100001;
            15'd30245: log10_cal = 16'b0000010111100001;
            15'd30246: log10_cal = 16'b0000010111100001;
            15'd30247: log10_cal = 16'b0000010111100001;
            15'd30248: log10_cal = 16'b0000010111100001;
            15'd30249: log10_cal = 16'b0000010111100001;
            15'd30250: log10_cal = 16'b0000010111100001;
            15'd30251: log10_cal = 16'b0000010111100001;
            15'd30252: log10_cal = 16'b0000010111100001;
            15'd30253: log10_cal = 16'b0000010111100001;
            15'd30254: log10_cal = 16'b0000010111100001;
            15'd30255: log10_cal = 16'b0000010111100001;
            15'd30256: log10_cal = 16'b0000010111100001;
            15'd30257: log10_cal = 16'b0000010111100001;
            15'd30258: log10_cal = 16'b0000010111100001;
            15'd30259: log10_cal = 16'b0000010111100001;
            15'd30260: log10_cal = 16'b0000010111100001;
            15'd30261: log10_cal = 16'b0000010111100001;
            15'd30262: log10_cal = 16'b0000010111100001;
            15'd30263: log10_cal = 16'b0000010111100001;
            15'd30264: log10_cal = 16'b0000010111100001;
            15'd30265: log10_cal = 16'b0000010111100001;
            15'd30266: log10_cal = 16'b0000010111100001;
            15'd30267: log10_cal = 16'b0000010111100001;
            15'd30268: log10_cal = 16'b0000010111100001;
            15'd30269: log10_cal = 16'b0000010111100001;
            15'd30270: log10_cal = 16'b0000010111100010;
            15'd30271: log10_cal = 16'b0000010111100010;
            15'd30272: log10_cal = 16'b0000010111100010;
            15'd30273: log10_cal = 16'b0000010111100010;
            15'd30274: log10_cal = 16'b0000010111100010;
            15'd30275: log10_cal = 16'b0000010111100010;
            15'd30276: log10_cal = 16'b0000010111100010;
            15'd30277: log10_cal = 16'b0000010111100010;
            15'd30278: log10_cal = 16'b0000010111100010;
            15'd30279: log10_cal = 16'b0000010111100010;
            15'd30280: log10_cal = 16'b0000010111100010;
            15'd30281: log10_cal = 16'b0000010111100010;
            15'd30282: log10_cal = 16'b0000010111100010;
            15'd30283: log10_cal = 16'b0000010111100010;
            15'd30284: log10_cal = 16'b0000010111100010;
            15'd30285: log10_cal = 16'b0000010111100010;
            15'd30286: log10_cal = 16'b0000010111100010;
            15'd30287: log10_cal = 16'b0000010111100010;
            15'd30288: log10_cal = 16'b0000010111100010;
            15'd30289: log10_cal = 16'b0000010111100010;
            15'd30290: log10_cal = 16'b0000010111100010;
            15'd30291: log10_cal = 16'b0000010111100010;
            15'd30292: log10_cal = 16'b0000010111100010;
            15'd30293: log10_cal = 16'b0000010111100010;
            15'd30294: log10_cal = 16'b0000010111100010;
            15'd30295: log10_cal = 16'b0000010111100010;
            15'd30296: log10_cal = 16'b0000010111100010;
            15'd30297: log10_cal = 16'b0000010111100010;
            15'd30298: log10_cal = 16'b0000010111100010;
            15'd30299: log10_cal = 16'b0000010111100010;
            15'd30300: log10_cal = 16'b0000010111100010;
            15'd30301: log10_cal = 16'b0000010111100010;
            15'd30302: log10_cal = 16'b0000010111100010;
            15'd30303: log10_cal = 16'b0000010111100010;
            15'd30304: log10_cal = 16'b0000010111100010;
            15'd30305: log10_cal = 16'b0000010111100010;
            15'd30306: log10_cal = 16'b0000010111100010;
            15'd30307: log10_cal = 16'b0000010111100010;
            15'd30308: log10_cal = 16'b0000010111100010;
            15'd30309: log10_cal = 16'b0000010111100010;
            15'd30310: log10_cal = 16'b0000010111100010;
            15'd30311: log10_cal = 16'b0000010111100010;
            15'd30312: log10_cal = 16'b0000010111100010;
            15'd30313: log10_cal = 16'b0000010111100010;
            15'd30314: log10_cal = 16'b0000010111100010;
            15'd30315: log10_cal = 16'b0000010111100010;
            15'd30316: log10_cal = 16'b0000010111100010;
            15'd30317: log10_cal = 16'b0000010111100010;
            15'd30318: log10_cal = 16'b0000010111100010;
            15'd30319: log10_cal = 16'b0000010111100010;
            15'd30320: log10_cal = 16'b0000010111100010;
            15'd30321: log10_cal = 16'b0000010111100010;
            15'd30322: log10_cal = 16'b0000010111100010;
            15'd30323: log10_cal = 16'b0000010111100010;
            15'd30324: log10_cal = 16'b0000010111100010;
            15'd30325: log10_cal = 16'b0000010111100010;
            15'd30326: log10_cal = 16'b0000010111100010;
            15'd30327: log10_cal = 16'b0000010111100010;
            15'd30328: log10_cal = 16'b0000010111100010;
            15'd30329: log10_cal = 16'b0000010111100010;
            15'd30330: log10_cal = 16'b0000010111100010;
            15'd30331: log10_cal = 16'b0000010111100010;
            15'd30332: log10_cal = 16'b0000010111100010;
            15'd30333: log10_cal = 16'b0000010111100010;
            15'd30334: log10_cal = 16'b0000010111100010;
            15'd30335: log10_cal = 16'b0000010111100010;
            15'd30336: log10_cal = 16'b0000010111100010;
            15'd30337: log10_cal = 16'b0000010111100010;
            15'd30338: log10_cal = 16'b0000010111100011;
            15'd30339: log10_cal = 16'b0000010111100011;
            15'd30340: log10_cal = 16'b0000010111100011;
            15'd30341: log10_cal = 16'b0000010111100011;
            15'd30342: log10_cal = 16'b0000010111100011;
            15'd30343: log10_cal = 16'b0000010111100011;
            15'd30344: log10_cal = 16'b0000010111100011;
            15'd30345: log10_cal = 16'b0000010111100011;
            15'd30346: log10_cal = 16'b0000010111100011;
            15'd30347: log10_cal = 16'b0000010111100011;
            15'd30348: log10_cal = 16'b0000010111100011;
            15'd30349: log10_cal = 16'b0000010111100011;
            15'd30350: log10_cal = 16'b0000010111100011;
            15'd30351: log10_cal = 16'b0000010111100011;
            15'd30352: log10_cal = 16'b0000010111100011;
            15'd30353: log10_cal = 16'b0000010111100011;
            15'd30354: log10_cal = 16'b0000010111100011;
            15'd30355: log10_cal = 16'b0000010111100011;
            15'd30356: log10_cal = 16'b0000010111100011;
            15'd30357: log10_cal = 16'b0000010111100011;
            15'd30358: log10_cal = 16'b0000010111100011;
            15'd30359: log10_cal = 16'b0000010111100011;
            15'd30360: log10_cal = 16'b0000010111100011;
            15'd30361: log10_cal = 16'b0000010111100011;
            15'd30362: log10_cal = 16'b0000010111100011;
            15'd30363: log10_cal = 16'b0000010111100011;
            15'd30364: log10_cal = 16'b0000010111100011;
            15'd30365: log10_cal = 16'b0000010111100011;
            15'd30366: log10_cal = 16'b0000010111100011;
            15'd30367: log10_cal = 16'b0000010111100011;
            15'd30368: log10_cal = 16'b0000010111100011;
            15'd30369: log10_cal = 16'b0000010111100011;
            15'd30370: log10_cal = 16'b0000010111100011;
            15'd30371: log10_cal = 16'b0000010111100011;
            15'd30372: log10_cal = 16'b0000010111100011;
            15'd30373: log10_cal = 16'b0000010111100011;
            15'd30374: log10_cal = 16'b0000010111100011;
            15'd30375: log10_cal = 16'b0000010111100011;
            15'd30376: log10_cal = 16'b0000010111100011;
            15'd30377: log10_cal = 16'b0000010111100011;
            15'd30378: log10_cal = 16'b0000010111100011;
            15'd30379: log10_cal = 16'b0000010111100011;
            15'd30380: log10_cal = 16'b0000010111100011;
            15'd30381: log10_cal = 16'b0000010111100011;
            15'd30382: log10_cal = 16'b0000010111100011;
            15'd30383: log10_cal = 16'b0000010111100011;
            15'd30384: log10_cal = 16'b0000010111100011;
            15'd30385: log10_cal = 16'b0000010111100011;
            15'd30386: log10_cal = 16'b0000010111100011;
            15'd30387: log10_cal = 16'b0000010111100011;
            15'd30388: log10_cal = 16'b0000010111100011;
            15'd30389: log10_cal = 16'b0000010111100011;
            15'd30390: log10_cal = 16'b0000010111100011;
            15'd30391: log10_cal = 16'b0000010111100011;
            15'd30392: log10_cal = 16'b0000010111100011;
            15'd30393: log10_cal = 16'b0000010111100011;
            15'd30394: log10_cal = 16'b0000010111100011;
            15'd30395: log10_cal = 16'b0000010111100011;
            15'd30396: log10_cal = 16'b0000010111100011;
            15'd30397: log10_cal = 16'b0000010111100011;
            15'd30398: log10_cal = 16'b0000010111100011;
            15'd30399: log10_cal = 16'b0000010111100011;
            15'd30400: log10_cal = 16'b0000010111100011;
            15'd30401: log10_cal = 16'b0000010111100011;
            15'd30402: log10_cal = 16'b0000010111100011;
            15'd30403: log10_cal = 16'b0000010111100011;
            15'd30404: log10_cal = 16'b0000010111100011;
            15'd30405: log10_cal = 16'b0000010111100011;
            15'd30406: log10_cal = 16'b0000010111100100;
            15'd30407: log10_cal = 16'b0000010111100100;
            15'd30408: log10_cal = 16'b0000010111100100;
            15'd30409: log10_cal = 16'b0000010111100100;
            15'd30410: log10_cal = 16'b0000010111100100;
            15'd30411: log10_cal = 16'b0000010111100100;
            15'd30412: log10_cal = 16'b0000010111100100;
            15'd30413: log10_cal = 16'b0000010111100100;
            15'd30414: log10_cal = 16'b0000010111100100;
            15'd30415: log10_cal = 16'b0000010111100100;
            15'd30416: log10_cal = 16'b0000010111100100;
            15'd30417: log10_cal = 16'b0000010111100100;
            15'd30418: log10_cal = 16'b0000010111100100;
            15'd30419: log10_cal = 16'b0000010111100100;
            15'd30420: log10_cal = 16'b0000010111100100;
            15'd30421: log10_cal = 16'b0000010111100100;
            15'd30422: log10_cal = 16'b0000010111100100;
            15'd30423: log10_cal = 16'b0000010111100100;
            15'd30424: log10_cal = 16'b0000010111100100;
            15'd30425: log10_cal = 16'b0000010111100100;
            15'd30426: log10_cal = 16'b0000010111100100;
            15'd30427: log10_cal = 16'b0000010111100100;
            15'd30428: log10_cal = 16'b0000010111100100;
            15'd30429: log10_cal = 16'b0000010111100100;
            15'd30430: log10_cal = 16'b0000010111100100;
            15'd30431: log10_cal = 16'b0000010111100100;
            15'd30432: log10_cal = 16'b0000010111100100;
            15'd30433: log10_cal = 16'b0000010111100100;
            15'd30434: log10_cal = 16'b0000010111100100;
            15'd30435: log10_cal = 16'b0000010111100100;
            15'd30436: log10_cal = 16'b0000010111100100;
            15'd30437: log10_cal = 16'b0000010111100100;
            15'd30438: log10_cal = 16'b0000010111100100;
            15'd30439: log10_cal = 16'b0000010111100100;
            15'd30440: log10_cal = 16'b0000010111100100;
            15'd30441: log10_cal = 16'b0000010111100100;
            15'd30442: log10_cal = 16'b0000010111100100;
            15'd30443: log10_cal = 16'b0000010111100100;
            15'd30444: log10_cal = 16'b0000010111100100;
            15'd30445: log10_cal = 16'b0000010111100100;
            15'd30446: log10_cal = 16'b0000010111100100;
            15'd30447: log10_cal = 16'b0000010111100100;
            15'd30448: log10_cal = 16'b0000010111100100;
            15'd30449: log10_cal = 16'b0000010111100100;
            15'd30450: log10_cal = 16'b0000010111100100;
            15'd30451: log10_cal = 16'b0000010111100100;
            15'd30452: log10_cal = 16'b0000010111100100;
            15'd30453: log10_cal = 16'b0000010111100100;
            15'd30454: log10_cal = 16'b0000010111100100;
            15'd30455: log10_cal = 16'b0000010111100100;
            15'd30456: log10_cal = 16'b0000010111100100;
            15'd30457: log10_cal = 16'b0000010111100100;
            15'd30458: log10_cal = 16'b0000010111100100;
            15'd30459: log10_cal = 16'b0000010111100100;
            15'd30460: log10_cal = 16'b0000010111100100;
            15'd30461: log10_cal = 16'b0000010111100100;
            15'd30462: log10_cal = 16'b0000010111100100;
            15'd30463: log10_cal = 16'b0000010111100100;
            15'd30464: log10_cal = 16'b0000010111100100;
            15'd30465: log10_cal = 16'b0000010111100100;
            15'd30466: log10_cal = 16'b0000010111100100;
            15'd30467: log10_cal = 16'b0000010111100100;
            15'd30468: log10_cal = 16'b0000010111100100;
            15'd30469: log10_cal = 16'b0000010111100100;
            15'd30470: log10_cal = 16'b0000010111100100;
            15'd30471: log10_cal = 16'b0000010111100100;
            15'd30472: log10_cal = 16'b0000010111100100;
            15'd30473: log10_cal = 16'b0000010111100100;
            15'd30474: log10_cal = 16'b0000010111100100;
            15'd30475: log10_cal = 16'b0000010111100101;
            15'd30476: log10_cal = 16'b0000010111100101;
            15'd30477: log10_cal = 16'b0000010111100101;
            15'd30478: log10_cal = 16'b0000010111100101;
            15'd30479: log10_cal = 16'b0000010111100101;
            15'd30480: log10_cal = 16'b0000010111100101;
            15'd30481: log10_cal = 16'b0000010111100101;
            15'd30482: log10_cal = 16'b0000010111100101;
            15'd30483: log10_cal = 16'b0000010111100101;
            15'd30484: log10_cal = 16'b0000010111100101;
            15'd30485: log10_cal = 16'b0000010111100101;
            15'd30486: log10_cal = 16'b0000010111100101;
            15'd30487: log10_cal = 16'b0000010111100101;
            15'd30488: log10_cal = 16'b0000010111100101;
            15'd30489: log10_cal = 16'b0000010111100101;
            15'd30490: log10_cal = 16'b0000010111100101;
            15'd30491: log10_cal = 16'b0000010111100101;
            15'd30492: log10_cal = 16'b0000010111100101;
            15'd30493: log10_cal = 16'b0000010111100101;
            15'd30494: log10_cal = 16'b0000010111100101;
            15'd30495: log10_cal = 16'b0000010111100101;
            15'd30496: log10_cal = 16'b0000010111100101;
            15'd30497: log10_cal = 16'b0000010111100101;
            15'd30498: log10_cal = 16'b0000010111100101;
            15'd30499: log10_cal = 16'b0000010111100101;
            15'd30500: log10_cal = 16'b0000010111100101;
            15'd30501: log10_cal = 16'b0000010111100101;
            15'd30502: log10_cal = 16'b0000010111100101;
            15'd30503: log10_cal = 16'b0000010111100101;
            15'd30504: log10_cal = 16'b0000010111100101;
            15'd30505: log10_cal = 16'b0000010111100101;
            15'd30506: log10_cal = 16'b0000010111100101;
            15'd30507: log10_cal = 16'b0000010111100101;
            15'd30508: log10_cal = 16'b0000010111100101;
            15'd30509: log10_cal = 16'b0000010111100101;
            15'd30510: log10_cal = 16'b0000010111100101;
            15'd30511: log10_cal = 16'b0000010111100101;
            15'd30512: log10_cal = 16'b0000010111100101;
            15'd30513: log10_cal = 16'b0000010111100101;
            15'd30514: log10_cal = 16'b0000010111100101;
            15'd30515: log10_cal = 16'b0000010111100101;
            15'd30516: log10_cal = 16'b0000010111100101;
            15'd30517: log10_cal = 16'b0000010111100101;
            15'd30518: log10_cal = 16'b0000010111100101;
            15'd30519: log10_cal = 16'b0000010111100101;
            15'd30520: log10_cal = 16'b0000010111100101;
            15'd30521: log10_cal = 16'b0000010111100101;
            15'd30522: log10_cal = 16'b0000010111100101;
            15'd30523: log10_cal = 16'b0000010111100101;
            15'd30524: log10_cal = 16'b0000010111100101;
            15'd30525: log10_cal = 16'b0000010111100101;
            15'd30526: log10_cal = 16'b0000010111100101;
            15'd30527: log10_cal = 16'b0000010111100101;
            15'd30528: log10_cal = 16'b0000010111100101;
            15'd30529: log10_cal = 16'b0000010111100101;
            15'd30530: log10_cal = 16'b0000010111100101;
            15'd30531: log10_cal = 16'b0000010111100101;
            15'd30532: log10_cal = 16'b0000010111100101;
            15'd30533: log10_cal = 16'b0000010111100101;
            15'd30534: log10_cal = 16'b0000010111100101;
            15'd30535: log10_cal = 16'b0000010111100101;
            15'd30536: log10_cal = 16'b0000010111100101;
            15'd30537: log10_cal = 16'b0000010111100101;
            15'd30538: log10_cal = 16'b0000010111100101;
            15'd30539: log10_cal = 16'b0000010111100101;
            15'd30540: log10_cal = 16'b0000010111100101;
            15'd30541: log10_cal = 16'b0000010111100101;
            15'd30542: log10_cal = 16'b0000010111100101;
            15'd30543: log10_cal = 16'b0000010111100110;
            15'd30544: log10_cal = 16'b0000010111100110;
            15'd30545: log10_cal = 16'b0000010111100110;
            15'd30546: log10_cal = 16'b0000010111100110;
            15'd30547: log10_cal = 16'b0000010111100110;
            15'd30548: log10_cal = 16'b0000010111100110;
            15'd30549: log10_cal = 16'b0000010111100110;
            15'd30550: log10_cal = 16'b0000010111100110;
            15'd30551: log10_cal = 16'b0000010111100110;
            15'd30552: log10_cal = 16'b0000010111100110;
            15'd30553: log10_cal = 16'b0000010111100110;
            15'd30554: log10_cal = 16'b0000010111100110;
            15'd30555: log10_cal = 16'b0000010111100110;
            15'd30556: log10_cal = 16'b0000010111100110;
            15'd30557: log10_cal = 16'b0000010111100110;
            15'd30558: log10_cal = 16'b0000010111100110;
            15'd30559: log10_cal = 16'b0000010111100110;
            15'd30560: log10_cal = 16'b0000010111100110;
            15'd30561: log10_cal = 16'b0000010111100110;
            15'd30562: log10_cal = 16'b0000010111100110;
            15'd30563: log10_cal = 16'b0000010111100110;
            15'd30564: log10_cal = 16'b0000010111100110;
            15'd30565: log10_cal = 16'b0000010111100110;
            15'd30566: log10_cal = 16'b0000010111100110;
            15'd30567: log10_cal = 16'b0000010111100110;
            15'd30568: log10_cal = 16'b0000010111100110;
            15'd30569: log10_cal = 16'b0000010111100110;
            15'd30570: log10_cal = 16'b0000010111100110;
            15'd30571: log10_cal = 16'b0000010111100110;
            15'd30572: log10_cal = 16'b0000010111100110;
            15'd30573: log10_cal = 16'b0000010111100110;
            15'd30574: log10_cal = 16'b0000010111100110;
            15'd30575: log10_cal = 16'b0000010111100110;
            15'd30576: log10_cal = 16'b0000010111100110;
            15'd30577: log10_cal = 16'b0000010111100110;
            15'd30578: log10_cal = 16'b0000010111100110;
            15'd30579: log10_cal = 16'b0000010111100110;
            15'd30580: log10_cal = 16'b0000010111100110;
            15'd30581: log10_cal = 16'b0000010111100110;
            15'd30582: log10_cal = 16'b0000010111100110;
            15'd30583: log10_cal = 16'b0000010111100110;
            15'd30584: log10_cal = 16'b0000010111100110;
            15'd30585: log10_cal = 16'b0000010111100110;
            15'd30586: log10_cal = 16'b0000010111100110;
            15'd30587: log10_cal = 16'b0000010111100110;
            15'd30588: log10_cal = 16'b0000010111100110;
            15'd30589: log10_cal = 16'b0000010111100110;
            15'd30590: log10_cal = 16'b0000010111100110;
            15'd30591: log10_cal = 16'b0000010111100110;
            15'd30592: log10_cal = 16'b0000010111100110;
            15'd30593: log10_cal = 16'b0000010111100110;
            15'd30594: log10_cal = 16'b0000010111100110;
            15'd30595: log10_cal = 16'b0000010111100110;
            15'd30596: log10_cal = 16'b0000010111100110;
            15'd30597: log10_cal = 16'b0000010111100110;
            15'd30598: log10_cal = 16'b0000010111100110;
            15'd30599: log10_cal = 16'b0000010111100110;
            15'd30600: log10_cal = 16'b0000010111100110;
            15'd30601: log10_cal = 16'b0000010111100110;
            15'd30602: log10_cal = 16'b0000010111100110;
            15'd30603: log10_cal = 16'b0000010111100110;
            15'd30604: log10_cal = 16'b0000010111100110;
            15'd30605: log10_cal = 16'b0000010111100110;
            15'd30606: log10_cal = 16'b0000010111100110;
            15'd30607: log10_cal = 16'b0000010111100110;
            15'd30608: log10_cal = 16'b0000010111100110;
            15'd30609: log10_cal = 16'b0000010111100110;
            15'd30610: log10_cal = 16'b0000010111100110;
            15'd30611: log10_cal = 16'b0000010111100110;
            15'd30612: log10_cal = 16'b0000010111100111;
            15'd30613: log10_cal = 16'b0000010111100111;
            15'd30614: log10_cal = 16'b0000010111100111;
            15'd30615: log10_cal = 16'b0000010111100111;
            15'd30616: log10_cal = 16'b0000010111100111;
            15'd30617: log10_cal = 16'b0000010111100111;
            15'd30618: log10_cal = 16'b0000010111100111;
            15'd30619: log10_cal = 16'b0000010111100111;
            15'd30620: log10_cal = 16'b0000010111100111;
            15'd30621: log10_cal = 16'b0000010111100111;
            15'd30622: log10_cal = 16'b0000010111100111;
            15'd30623: log10_cal = 16'b0000010111100111;
            15'd30624: log10_cal = 16'b0000010111100111;
            15'd30625: log10_cal = 16'b0000010111100111;
            15'd30626: log10_cal = 16'b0000010111100111;
            15'd30627: log10_cal = 16'b0000010111100111;
            15'd30628: log10_cal = 16'b0000010111100111;
            15'd30629: log10_cal = 16'b0000010111100111;
            15'd30630: log10_cal = 16'b0000010111100111;
            15'd30631: log10_cal = 16'b0000010111100111;
            15'd30632: log10_cal = 16'b0000010111100111;
            15'd30633: log10_cal = 16'b0000010111100111;
            15'd30634: log10_cal = 16'b0000010111100111;
            15'd30635: log10_cal = 16'b0000010111100111;
            15'd30636: log10_cal = 16'b0000010111100111;
            15'd30637: log10_cal = 16'b0000010111100111;
            15'd30638: log10_cal = 16'b0000010111100111;
            15'd30639: log10_cal = 16'b0000010111100111;
            15'd30640: log10_cal = 16'b0000010111100111;
            15'd30641: log10_cal = 16'b0000010111100111;
            15'd30642: log10_cal = 16'b0000010111100111;
            15'd30643: log10_cal = 16'b0000010111100111;
            15'd30644: log10_cal = 16'b0000010111100111;
            15'd30645: log10_cal = 16'b0000010111100111;
            15'd30646: log10_cal = 16'b0000010111100111;
            15'd30647: log10_cal = 16'b0000010111100111;
            15'd30648: log10_cal = 16'b0000010111100111;
            15'd30649: log10_cal = 16'b0000010111100111;
            15'd30650: log10_cal = 16'b0000010111100111;
            15'd30651: log10_cal = 16'b0000010111100111;
            15'd30652: log10_cal = 16'b0000010111100111;
            15'd30653: log10_cal = 16'b0000010111100111;
            15'd30654: log10_cal = 16'b0000010111100111;
            15'd30655: log10_cal = 16'b0000010111100111;
            15'd30656: log10_cal = 16'b0000010111100111;
            15'd30657: log10_cal = 16'b0000010111100111;
            15'd30658: log10_cal = 16'b0000010111100111;
            15'd30659: log10_cal = 16'b0000010111100111;
            15'd30660: log10_cal = 16'b0000010111100111;
            15'd30661: log10_cal = 16'b0000010111100111;
            15'd30662: log10_cal = 16'b0000010111100111;
            15'd30663: log10_cal = 16'b0000010111100111;
            15'd30664: log10_cal = 16'b0000010111100111;
            15'd30665: log10_cal = 16'b0000010111100111;
            15'd30666: log10_cal = 16'b0000010111100111;
            15'd30667: log10_cal = 16'b0000010111100111;
            15'd30668: log10_cal = 16'b0000010111100111;
            15'd30669: log10_cal = 16'b0000010111100111;
            15'd30670: log10_cal = 16'b0000010111100111;
            15'd30671: log10_cal = 16'b0000010111100111;
            15'd30672: log10_cal = 16'b0000010111100111;
            15'd30673: log10_cal = 16'b0000010111100111;
            15'd30674: log10_cal = 16'b0000010111100111;
            15'd30675: log10_cal = 16'b0000010111100111;
            15'd30676: log10_cal = 16'b0000010111100111;
            15'd30677: log10_cal = 16'b0000010111100111;
            15'd30678: log10_cal = 16'b0000010111100111;
            15'd30679: log10_cal = 16'b0000010111100111;
            15'd30680: log10_cal = 16'b0000010111100111;
            15'd30681: log10_cal = 16'b0000010111101000;
            15'd30682: log10_cal = 16'b0000010111101000;
            15'd30683: log10_cal = 16'b0000010111101000;
            15'd30684: log10_cal = 16'b0000010111101000;
            15'd30685: log10_cal = 16'b0000010111101000;
            15'd30686: log10_cal = 16'b0000010111101000;
            15'd30687: log10_cal = 16'b0000010111101000;
            15'd30688: log10_cal = 16'b0000010111101000;
            15'd30689: log10_cal = 16'b0000010111101000;
            15'd30690: log10_cal = 16'b0000010111101000;
            15'd30691: log10_cal = 16'b0000010111101000;
            15'd30692: log10_cal = 16'b0000010111101000;
            15'd30693: log10_cal = 16'b0000010111101000;
            15'd30694: log10_cal = 16'b0000010111101000;
            15'd30695: log10_cal = 16'b0000010111101000;
            15'd30696: log10_cal = 16'b0000010111101000;
            15'd30697: log10_cal = 16'b0000010111101000;
            15'd30698: log10_cal = 16'b0000010111101000;
            15'd30699: log10_cal = 16'b0000010111101000;
            15'd30700: log10_cal = 16'b0000010111101000;
            15'd30701: log10_cal = 16'b0000010111101000;
            15'd30702: log10_cal = 16'b0000010111101000;
            15'd30703: log10_cal = 16'b0000010111101000;
            15'd30704: log10_cal = 16'b0000010111101000;
            15'd30705: log10_cal = 16'b0000010111101000;
            15'd30706: log10_cal = 16'b0000010111101000;
            15'd30707: log10_cal = 16'b0000010111101000;
            15'd30708: log10_cal = 16'b0000010111101000;
            15'd30709: log10_cal = 16'b0000010111101000;
            15'd30710: log10_cal = 16'b0000010111101000;
            15'd30711: log10_cal = 16'b0000010111101000;
            15'd30712: log10_cal = 16'b0000010111101000;
            15'd30713: log10_cal = 16'b0000010111101000;
            15'd30714: log10_cal = 16'b0000010111101000;
            15'd30715: log10_cal = 16'b0000010111101000;
            15'd30716: log10_cal = 16'b0000010111101000;
            15'd30717: log10_cal = 16'b0000010111101000;
            15'd30718: log10_cal = 16'b0000010111101000;
            15'd30719: log10_cal = 16'b0000010111101000;
            15'd30720: log10_cal = 16'b0000010111101000;
            15'd30721: log10_cal = 16'b0000010111101000;
            15'd30722: log10_cal = 16'b0000010111101000;
            15'd30723: log10_cal = 16'b0000010111101000;
            15'd30724: log10_cal = 16'b0000010111101000;
            15'd30725: log10_cal = 16'b0000010111101000;
            15'd30726: log10_cal = 16'b0000010111101000;
            15'd30727: log10_cal = 16'b0000010111101000;
            15'd30728: log10_cal = 16'b0000010111101000;
            15'd30729: log10_cal = 16'b0000010111101000;
            15'd30730: log10_cal = 16'b0000010111101000;
            15'd30731: log10_cal = 16'b0000010111101000;
            15'd30732: log10_cal = 16'b0000010111101000;
            15'd30733: log10_cal = 16'b0000010111101000;
            15'd30734: log10_cal = 16'b0000010111101000;
            15'd30735: log10_cal = 16'b0000010111101000;
            15'd30736: log10_cal = 16'b0000010111101000;
            15'd30737: log10_cal = 16'b0000010111101000;
            15'd30738: log10_cal = 16'b0000010111101000;
            15'd30739: log10_cal = 16'b0000010111101000;
            15'd30740: log10_cal = 16'b0000010111101000;
            15'd30741: log10_cal = 16'b0000010111101000;
            15'd30742: log10_cal = 16'b0000010111101000;
            15'd30743: log10_cal = 16'b0000010111101000;
            15'd30744: log10_cal = 16'b0000010111101000;
            15'd30745: log10_cal = 16'b0000010111101000;
            15'd30746: log10_cal = 16'b0000010111101000;
            15'd30747: log10_cal = 16'b0000010111101000;
            15'd30748: log10_cal = 16'b0000010111101000;
            15'd30749: log10_cal = 16'b0000010111101000;
            15'd30750: log10_cal = 16'b0000010111101001;
            15'd30751: log10_cal = 16'b0000010111101001;
            15'd30752: log10_cal = 16'b0000010111101001;
            15'd30753: log10_cal = 16'b0000010111101001;
            15'd30754: log10_cal = 16'b0000010111101001;
            15'd30755: log10_cal = 16'b0000010111101001;
            15'd30756: log10_cal = 16'b0000010111101001;
            15'd30757: log10_cal = 16'b0000010111101001;
            15'd30758: log10_cal = 16'b0000010111101001;
            15'd30759: log10_cal = 16'b0000010111101001;
            15'd30760: log10_cal = 16'b0000010111101001;
            15'd30761: log10_cal = 16'b0000010111101001;
            15'd30762: log10_cal = 16'b0000010111101001;
            15'd30763: log10_cal = 16'b0000010111101001;
            15'd30764: log10_cal = 16'b0000010111101001;
            15'd30765: log10_cal = 16'b0000010111101001;
            15'd30766: log10_cal = 16'b0000010111101001;
            15'd30767: log10_cal = 16'b0000010111101001;
            15'd30768: log10_cal = 16'b0000010111101001;
            15'd30769: log10_cal = 16'b0000010111101001;
            15'd30770: log10_cal = 16'b0000010111101001;
            15'd30771: log10_cal = 16'b0000010111101001;
            15'd30772: log10_cal = 16'b0000010111101001;
            15'd30773: log10_cal = 16'b0000010111101001;
            15'd30774: log10_cal = 16'b0000010111101001;
            15'd30775: log10_cal = 16'b0000010111101001;
            15'd30776: log10_cal = 16'b0000010111101001;
            15'd30777: log10_cal = 16'b0000010111101001;
            15'd30778: log10_cal = 16'b0000010111101001;
            15'd30779: log10_cal = 16'b0000010111101001;
            15'd30780: log10_cal = 16'b0000010111101001;
            15'd30781: log10_cal = 16'b0000010111101001;
            15'd30782: log10_cal = 16'b0000010111101001;
            15'd30783: log10_cal = 16'b0000010111101001;
            15'd30784: log10_cal = 16'b0000010111101001;
            15'd30785: log10_cal = 16'b0000010111101001;
            15'd30786: log10_cal = 16'b0000010111101001;
            15'd30787: log10_cal = 16'b0000010111101001;
            15'd30788: log10_cal = 16'b0000010111101001;
            15'd30789: log10_cal = 16'b0000010111101001;
            15'd30790: log10_cal = 16'b0000010111101001;
            15'd30791: log10_cal = 16'b0000010111101001;
            15'd30792: log10_cal = 16'b0000010111101001;
            15'd30793: log10_cal = 16'b0000010111101001;
            15'd30794: log10_cal = 16'b0000010111101001;
            15'd30795: log10_cal = 16'b0000010111101001;
            15'd30796: log10_cal = 16'b0000010111101001;
            15'd30797: log10_cal = 16'b0000010111101001;
            15'd30798: log10_cal = 16'b0000010111101001;
            15'd30799: log10_cal = 16'b0000010111101001;
            15'd30800: log10_cal = 16'b0000010111101001;
            15'd30801: log10_cal = 16'b0000010111101001;
            15'd30802: log10_cal = 16'b0000010111101001;
            15'd30803: log10_cal = 16'b0000010111101001;
            15'd30804: log10_cal = 16'b0000010111101001;
            15'd30805: log10_cal = 16'b0000010111101001;
            15'd30806: log10_cal = 16'b0000010111101001;
            15'd30807: log10_cal = 16'b0000010111101001;
            15'd30808: log10_cal = 16'b0000010111101001;
            15'd30809: log10_cal = 16'b0000010111101001;
            15'd30810: log10_cal = 16'b0000010111101001;
            15'd30811: log10_cal = 16'b0000010111101001;
            15'd30812: log10_cal = 16'b0000010111101001;
            15'd30813: log10_cal = 16'b0000010111101001;
            15'd30814: log10_cal = 16'b0000010111101001;
            15'd30815: log10_cal = 16'b0000010111101001;
            15'd30816: log10_cal = 16'b0000010111101001;
            15'd30817: log10_cal = 16'b0000010111101001;
            15'd30818: log10_cal = 16'b0000010111101001;
            15'd30819: log10_cal = 16'b0000010111101010;
            15'd30820: log10_cal = 16'b0000010111101010;
            15'd30821: log10_cal = 16'b0000010111101010;
            15'd30822: log10_cal = 16'b0000010111101010;
            15'd30823: log10_cal = 16'b0000010111101010;
            15'd30824: log10_cal = 16'b0000010111101010;
            15'd30825: log10_cal = 16'b0000010111101010;
            15'd30826: log10_cal = 16'b0000010111101010;
            15'd30827: log10_cal = 16'b0000010111101010;
            15'd30828: log10_cal = 16'b0000010111101010;
            15'd30829: log10_cal = 16'b0000010111101010;
            15'd30830: log10_cal = 16'b0000010111101010;
            15'd30831: log10_cal = 16'b0000010111101010;
            15'd30832: log10_cal = 16'b0000010111101010;
            15'd30833: log10_cal = 16'b0000010111101010;
            15'd30834: log10_cal = 16'b0000010111101010;
            15'd30835: log10_cal = 16'b0000010111101010;
            15'd30836: log10_cal = 16'b0000010111101010;
            15'd30837: log10_cal = 16'b0000010111101010;
            15'd30838: log10_cal = 16'b0000010111101010;
            15'd30839: log10_cal = 16'b0000010111101010;
            15'd30840: log10_cal = 16'b0000010111101010;
            15'd30841: log10_cal = 16'b0000010111101010;
            15'd30842: log10_cal = 16'b0000010111101010;
            15'd30843: log10_cal = 16'b0000010111101010;
            15'd30844: log10_cal = 16'b0000010111101010;
            15'd30845: log10_cal = 16'b0000010111101010;
            15'd30846: log10_cal = 16'b0000010111101010;
            15'd30847: log10_cal = 16'b0000010111101010;
            15'd30848: log10_cal = 16'b0000010111101010;
            15'd30849: log10_cal = 16'b0000010111101010;
            15'd30850: log10_cal = 16'b0000010111101010;
            15'd30851: log10_cal = 16'b0000010111101010;
            15'd30852: log10_cal = 16'b0000010111101010;
            15'd30853: log10_cal = 16'b0000010111101010;
            15'd30854: log10_cal = 16'b0000010111101010;
            15'd30855: log10_cal = 16'b0000010111101010;
            15'd30856: log10_cal = 16'b0000010111101010;
            15'd30857: log10_cal = 16'b0000010111101010;
            15'd30858: log10_cal = 16'b0000010111101010;
            15'd30859: log10_cal = 16'b0000010111101010;
            15'd30860: log10_cal = 16'b0000010111101010;
            15'd30861: log10_cal = 16'b0000010111101010;
            15'd30862: log10_cal = 16'b0000010111101010;
            15'd30863: log10_cal = 16'b0000010111101010;
            15'd30864: log10_cal = 16'b0000010111101010;
            15'd30865: log10_cal = 16'b0000010111101010;
            15'd30866: log10_cal = 16'b0000010111101010;
            15'd30867: log10_cal = 16'b0000010111101010;
            15'd30868: log10_cal = 16'b0000010111101010;
            15'd30869: log10_cal = 16'b0000010111101010;
            15'd30870: log10_cal = 16'b0000010111101010;
            15'd30871: log10_cal = 16'b0000010111101010;
            15'd30872: log10_cal = 16'b0000010111101010;
            15'd30873: log10_cal = 16'b0000010111101010;
            15'd30874: log10_cal = 16'b0000010111101010;
            15'd30875: log10_cal = 16'b0000010111101010;
            15'd30876: log10_cal = 16'b0000010111101010;
            15'd30877: log10_cal = 16'b0000010111101010;
            15'd30878: log10_cal = 16'b0000010111101010;
            15'd30879: log10_cal = 16'b0000010111101010;
            15'd30880: log10_cal = 16'b0000010111101010;
            15'd30881: log10_cal = 16'b0000010111101010;
            15'd30882: log10_cal = 16'b0000010111101010;
            15'd30883: log10_cal = 16'b0000010111101010;
            15'd30884: log10_cal = 16'b0000010111101010;
            15'd30885: log10_cal = 16'b0000010111101010;
            15'd30886: log10_cal = 16'b0000010111101010;
            15'd30887: log10_cal = 16'b0000010111101010;
            15'd30888: log10_cal = 16'b0000010111101010;
            15'd30889: log10_cal = 16'b0000010111101011;
            15'd30890: log10_cal = 16'b0000010111101011;
            15'd30891: log10_cal = 16'b0000010111101011;
            15'd30892: log10_cal = 16'b0000010111101011;
            15'd30893: log10_cal = 16'b0000010111101011;
            15'd30894: log10_cal = 16'b0000010111101011;
            15'd30895: log10_cal = 16'b0000010111101011;
            15'd30896: log10_cal = 16'b0000010111101011;
            15'd30897: log10_cal = 16'b0000010111101011;
            15'd30898: log10_cal = 16'b0000010111101011;
            15'd30899: log10_cal = 16'b0000010111101011;
            15'd30900: log10_cal = 16'b0000010111101011;
            15'd30901: log10_cal = 16'b0000010111101011;
            15'd30902: log10_cal = 16'b0000010111101011;
            15'd30903: log10_cal = 16'b0000010111101011;
            15'd30904: log10_cal = 16'b0000010111101011;
            15'd30905: log10_cal = 16'b0000010111101011;
            15'd30906: log10_cal = 16'b0000010111101011;
            15'd30907: log10_cal = 16'b0000010111101011;
            15'd30908: log10_cal = 16'b0000010111101011;
            15'd30909: log10_cal = 16'b0000010111101011;
            15'd30910: log10_cal = 16'b0000010111101011;
            15'd30911: log10_cal = 16'b0000010111101011;
            15'd30912: log10_cal = 16'b0000010111101011;
            15'd30913: log10_cal = 16'b0000010111101011;
            15'd30914: log10_cal = 16'b0000010111101011;
            15'd30915: log10_cal = 16'b0000010111101011;
            15'd30916: log10_cal = 16'b0000010111101011;
            15'd30917: log10_cal = 16'b0000010111101011;
            15'd30918: log10_cal = 16'b0000010111101011;
            15'd30919: log10_cal = 16'b0000010111101011;
            15'd30920: log10_cal = 16'b0000010111101011;
            15'd30921: log10_cal = 16'b0000010111101011;
            15'd30922: log10_cal = 16'b0000010111101011;
            15'd30923: log10_cal = 16'b0000010111101011;
            15'd30924: log10_cal = 16'b0000010111101011;
            15'd30925: log10_cal = 16'b0000010111101011;
            15'd30926: log10_cal = 16'b0000010111101011;
            15'd30927: log10_cal = 16'b0000010111101011;
            15'd30928: log10_cal = 16'b0000010111101011;
            15'd30929: log10_cal = 16'b0000010111101011;
            15'd30930: log10_cal = 16'b0000010111101011;
            15'd30931: log10_cal = 16'b0000010111101011;
            15'd30932: log10_cal = 16'b0000010111101011;
            15'd30933: log10_cal = 16'b0000010111101011;
            15'd30934: log10_cal = 16'b0000010111101011;
            15'd30935: log10_cal = 16'b0000010111101011;
            15'd30936: log10_cal = 16'b0000010111101011;
            15'd30937: log10_cal = 16'b0000010111101011;
            15'd30938: log10_cal = 16'b0000010111101011;
            15'd30939: log10_cal = 16'b0000010111101011;
            15'd30940: log10_cal = 16'b0000010111101011;
            15'd30941: log10_cal = 16'b0000010111101011;
            15'd30942: log10_cal = 16'b0000010111101011;
            15'd30943: log10_cal = 16'b0000010111101011;
            15'd30944: log10_cal = 16'b0000010111101011;
            15'd30945: log10_cal = 16'b0000010111101011;
            15'd30946: log10_cal = 16'b0000010111101011;
            15'd30947: log10_cal = 16'b0000010111101011;
            15'd30948: log10_cal = 16'b0000010111101011;
            15'd30949: log10_cal = 16'b0000010111101011;
            15'd30950: log10_cal = 16'b0000010111101011;
            15'd30951: log10_cal = 16'b0000010111101011;
            15'd30952: log10_cal = 16'b0000010111101011;
            15'd30953: log10_cal = 16'b0000010111101011;
            15'd30954: log10_cal = 16'b0000010111101011;
            15'd30955: log10_cal = 16'b0000010111101011;
            15'd30956: log10_cal = 16'b0000010111101011;
            15'd30957: log10_cal = 16'b0000010111101011;
            15'd30958: log10_cal = 16'b0000010111101100;
            15'd30959: log10_cal = 16'b0000010111101100;
            15'd30960: log10_cal = 16'b0000010111101100;
            15'd30961: log10_cal = 16'b0000010111101100;
            15'd30962: log10_cal = 16'b0000010111101100;
            15'd30963: log10_cal = 16'b0000010111101100;
            15'd30964: log10_cal = 16'b0000010111101100;
            15'd30965: log10_cal = 16'b0000010111101100;
            15'd30966: log10_cal = 16'b0000010111101100;
            15'd30967: log10_cal = 16'b0000010111101100;
            15'd30968: log10_cal = 16'b0000010111101100;
            15'd30969: log10_cal = 16'b0000010111101100;
            15'd30970: log10_cal = 16'b0000010111101100;
            15'd30971: log10_cal = 16'b0000010111101100;
            15'd30972: log10_cal = 16'b0000010111101100;
            15'd30973: log10_cal = 16'b0000010111101100;
            15'd30974: log10_cal = 16'b0000010111101100;
            15'd30975: log10_cal = 16'b0000010111101100;
            15'd30976: log10_cal = 16'b0000010111101100;
            15'd30977: log10_cal = 16'b0000010111101100;
            15'd30978: log10_cal = 16'b0000010111101100;
            15'd30979: log10_cal = 16'b0000010111101100;
            15'd30980: log10_cal = 16'b0000010111101100;
            15'd30981: log10_cal = 16'b0000010111101100;
            15'd30982: log10_cal = 16'b0000010111101100;
            15'd30983: log10_cal = 16'b0000010111101100;
            15'd30984: log10_cal = 16'b0000010111101100;
            15'd30985: log10_cal = 16'b0000010111101100;
            15'd30986: log10_cal = 16'b0000010111101100;
            15'd30987: log10_cal = 16'b0000010111101100;
            15'd30988: log10_cal = 16'b0000010111101100;
            15'd30989: log10_cal = 16'b0000010111101100;
            15'd30990: log10_cal = 16'b0000010111101100;
            15'd30991: log10_cal = 16'b0000010111101100;
            15'd30992: log10_cal = 16'b0000010111101100;
            15'd30993: log10_cal = 16'b0000010111101100;
            15'd30994: log10_cal = 16'b0000010111101100;
            15'd30995: log10_cal = 16'b0000010111101100;
            15'd30996: log10_cal = 16'b0000010111101100;
            15'd30997: log10_cal = 16'b0000010111101100;
            15'd30998: log10_cal = 16'b0000010111101100;
            15'd30999: log10_cal = 16'b0000010111101100;
            15'd31000: log10_cal = 16'b0000010111101100;
            15'd31001: log10_cal = 16'b0000010111101100;
            15'd31002: log10_cal = 16'b0000010111101100;
            15'd31003: log10_cal = 16'b0000010111101100;
            15'd31004: log10_cal = 16'b0000010111101100;
            15'd31005: log10_cal = 16'b0000010111101100;
            15'd31006: log10_cal = 16'b0000010111101100;
            15'd31007: log10_cal = 16'b0000010111101100;
            15'd31008: log10_cal = 16'b0000010111101100;
            15'd31009: log10_cal = 16'b0000010111101100;
            15'd31010: log10_cal = 16'b0000010111101100;
            15'd31011: log10_cal = 16'b0000010111101100;
            15'd31012: log10_cal = 16'b0000010111101100;
            15'd31013: log10_cal = 16'b0000010111101100;
            15'd31014: log10_cal = 16'b0000010111101100;
            15'd31015: log10_cal = 16'b0000010111101100;
            15'd31016: log10_cal = 16'b0000010111101100;
            15'd31017: log10_cal = 16'b0000010111101100;
            15'd31018: log10_cal = 16'b0000010111101100;
            15'd31019: log10_cal = 16'b0000010111101100;
            15'd31020: log10_cal = 16'b0000010111101100;
            15'd31021: log10_cal = 16'b0000010111101100;
            15'd31022: log10_cal = 16'b0000010111101100;
            15'd31023: log10_cal = 16'b0000010111101100;
            15'd31024: log10_cal = 16'b0000010111101100;
            15'd31025: log10_cal = 16'b0000010111101100;
            15'd31026: log10_cal = 16'b0000010111101100;
            15'd31027: log10_cal = 16'b0000010111101100;
            15'd31028: log10_cal = 16'b0000010111101101;
            15'd31029: log10_cal = 16'b0000010111101101;
            15'd31030: log10_cal = 16'b0000010111101101;
            15'd31031: log10_cal = 16'b0000010111101101;
            15'd31032: log10_cal = 16'b0000010111101101;
            15'd31033: log10_cal = 16'b0000010111101101;
            15'd31034: log10_cal = 16'b0000010111101101;
            15'd31035: log10_cal = 16'b0000010111101101;
            15'd31036: log10_cal = 16'b0000010111101101;
            15'd31037: log10_cal = 16'b0000010111101101;
            15'd31038: log10_cal = 16'b0000010111101101;
            15'd31039: log10_cal = 16'b0000010111101101;
            15'd31040: log10_cal = 16'b0000010111101101;
            15'd31041: log10_cal = 16'b0000010111101101;
            15'd31042: log10_cal = 16'b0000010111101101;
            15'd31043: log10_cal = 16'b0000010111101101;
            15'd31044: log10_cal = 16'b0000010111101101;
            15'd31045: log10_cal = 16'b0000010111101101;
            15'd31046: log10_cal = 16'b0000010111101101;
            15'd31047: log10_cal = 16'b0000010111101101;
            15'd31048: log10_cal = 16'b0000010111101101;
            15'd31049: log10_cal = 16'b0000010111101101;
            15'd31050: log10_cal = 16'b0000010111101101;
            15'd31051: log10_cal = 16'b0000010111101101;
            15'd31052: log10_cal = 16'b0000010111101101;
            15'd31053: log10_cal = 16'b0000010111101101;
            15'd31054: log10_cal = 16'b0000010111101101;
            15'd31055: log10_cal = 16'b0000010111101101;
            15'd31056: log10_cal = 16'b0000010111101101;
            15'd31057: log10_cal = 16'b0000010111101101;
            15'd31058: log10_cal = 16'b0000010111101101;
            15'd31059: log10_cal = 16'b0000010111101101;
            15'd31060: log10_cal = 16'b0000010111101101;
            15'd31061: log10_cal = 16'b0000010111101101;
            15'd31062: log10_cal = 16'b0000010111101101;
            15'd31063: log10_cal = 16'b0000010111101101;
            15'd31064: log10_cal = 16'b0000010111101101;
            15'd31065: log10_cal = 16'b0000010111101101;
            15'd31066: log10_cal = 16'b0000010111101101;
            15'd31067: log10_cal = 16'b0000010111101101;
            15'd31068: log10_cal = 16'b0000010111101101;
            15'd31069: log10_cal = 16'b0000010111101101;
            15'd31070: log10_cal = 16'b0000010111101101;
            15'd31071: log10_cal = 16'b0000010111101101;
            15'd31072: log10_cal = 16'b0000010111101101;
            15'd31073: log10_cal = 16'b0000010111101101;
            15'd31074: log10_cal = 16'b0000010111101101;
            15'd31075: log10_cal = 16'b0000010111101101;
            15'd31076: log10_cal = 16'b0000010111101101;
            15'd31077: log10_cal = 16'b0000010111101101;
            15'd31078: log10_cal = 16'b0000010111101101;
            15'd31079: log10_cal = 16'b0000010111101101;
            15'd31080: log10_cal = 16'b0000010111101101;
            15'd31081: log10_cal = 16'b0000010111101101;
            15'd31082: log10_cal = 16'b0000010111101101;
            15'd31083: log10_cal = 16'b0000010111101101;
            15'd31084: log10_cal = 16'b0000010111101101;
            15'd31085: log10_cal = 16'b0000010111101101;
            15'd31086: log10_cal = 16'b0000010111101101;
            15'd31087: log10_cal = 16'b0000010111101101;
            15'd31088: log10_cal = 16'b0000010111101101;
            15'd31089: log10_cal = 16'b0000010111101101;
            15'd31090: log10_cal = 16'b0000010111101101;
            15'd31091: log10_cal = 16'b0000010111101101;
            15'd31092: log10_cal = 16'b0000010111101101;
            15'd31093: log10_cal = 16'b0000010111101101;
            15'd31094: log10_cal = 16'b0000010111101101;
            15'd31095: log10_cal = 16'b0000010111101101;
            15'd31096: log10_cal = 16'b0000010111101101;
            15'd31097: log10_cal = 16'b0000010111101101;
            15'd31098: log10_cal = 16'b0000010111101110;
            15'd31099: log10_cal = 16'b0000010111101110;
            15'd31100: log10_cal = 16'b0000010111101110;
            15'd31101: log10_cal = 16'b0000010111101110;
            15'd31102: log10_cal = 16'b0000010111101110;
            15'd31103: log10_cal = 16'b0000010111101110;
            15'd31104: log10_cal = 16'b0000010111101110;
            15'd31105: log10_cal = 16'b0000010111101110;
            15'd31106: log10_cal = 16'b0000010111101110;
            15'd31107: log10_cal = 16'b0000010111101110;
            15'd31108: log10_cal = 16'b0000010111101110;
            15'd31109: log10_cal = 16'b0000010111101110;
            15'd31110: log10_cal = 16'b0000010111101110;
            15'd31111: log10_cal = 16'b0000010111101110;
            15'd31112: log10_cal = 16'b0000010111101110;
            15'd31113: log10_cal = 16'b0000010111101110;
            15'd31114: log10_cal = 16'b0000010111101110;
            15'd31115: log10_cal = 16'b0000010111101110;
            15'd31116: log10_cal = 16'b0000010111101110;
            15'd31117: log10_cal = 16'b0000010111101110;
            15'd31118: log10_cal = 16'b0000010111101110;
            15'd31119: log10_cal = 16'b0000010111101110;
            15'd31120: log10_cal = 16'b0000010111101110;
            15'd31121: log10_cal = 16'b0000010111101110;
            15'd31122: log10_cal = 16'b0000010111101110;
            15'd31123: log10_cal = 16'b0000010111101110;
            15'd31124: log10_cal = 16'b0000010111101110;
            15'd31125: log10_cal = 16'b0000010111101110;
            15'd31126: log10_cal = 16'b0000010111101110;
            15'd31127: log10_cal = 16'b0000010111101110;
            15'd31128: log10_cal = 16'b0000010111101110;
            15'd31129: log10_cal = 16'b0000010111101110;
            15'd31130: log10_cal = 16'b0000010111101110;
            15'd31131: log10_cal = 16'b0000010111101110;
            15'd31132: log10_cal = 16'b0000010111101110;
            15'd31133: log10_cal = 16'b0000010111101110;
            15'd31134: log10_cal = 16'b0000010111101110;
            15'd31135: log10_cal = 16'b0000010111101110;
            15'd31136: log10_cal = 16'b0000010111101110;
            15'd31137: log10_cal = 16'b0000010111101110;
            15'd31138: log10_cal = 16'b0000010111101110;
            15'd31139: log10_cal = 16'b0000010111101110;
            15'd31140: log10_cal = 16'b0000010111101110;
            15'd31141: log10_cal = 16'b0000010111101110;
            15'd31142: log10_cal = 16'b0000010111101110;
            15'd31143: log10_cal = 16'b0000010111101110;
            15'd31144: log10_cal = 16'b0000010111101110;
            15'd31145: log10_cal = 16'b0000010111101110;
            15'd31146: log10_cal = 16'b0000010111101110;
            15'd31147: log10_cal = 16'b0000010111101110;
            15'd31148: log10_cal = 16'b0000010111101110;
            15'd31149: log10_cal = 16'b0000010111101110;
            15'd31150: log10_cal = 16'b0000010111101110;
            15'd31151: log10_cal = 16'b0000010111101110;
            15'd31152: log10_cal = 16'b0000010111101110;
            15'd31153: log10_cal = 16'b0000010111101110;
            15'd31154: log10_cal = 16'b0000010111101110;
            15'd31155: log10_cal = 16'b0000010111101110;
            15'd31156: log10_cal = 16'b0000010111101110;
            15'd31157: log10_cal = 16'b0000010111101110;
            15'd31158: log10_cal = 16'b0000010111101110;
            15'd31159: log10_cal = 16'b0000010111101110;
            15'd31160: log10_cal = 16'b0000010111101110;
            15'd31161: log10_cal = 16'b0000010111101110;
            15'd31162: log10_cal = 16'b0000010111101110;
            15'd31163: log10_cal = 16'b0000010111101110;
            15'd31164: log10_cal = 16'b0000010111101110;
            15'd31165: log10_cal = 16'b0000010111101110;
            15'd31166: log10_cal = 16'b0000010111101110;
            15'd31167: log10_cal = 16'b0000010111101110;
            15'd31168: log10_cal = 16'b0000010111101111;
            15'd31169: log10_cal = 16'b0000010111101111;
            15'd31170: log10_cal = 16'b0000010111101111;
            15'd31171: log10_cal = 16'b0000010111101111;
            15'd31172: log10_cal = 16'b0000010111101111;
            15'd31173: log10_cal = 16'b0000010111101111;
            15'd31174: log10_cal = 16'b0000010111101111;
            15'd31175: log10_cal = 16'b0000010111101111;
            15'd31176: log10_cal = 16'b0000010111101111;
            15'd31177: log10_cal = 16'b0000010111101111;
            15'd31178: log10_cal = 16'b0000010111101111;
            15'd31179: log10_cal = 16'b0000010111101111;
            15'd31180: log10_cal = 16'b0000010111101111;
            15'd31181: log10_cal = 16'b0000010111101111;
            15'd31182: log10_cal = 16'b0000010111101111;
            15'd31183: log10_cal = 16'b0000010111101111;
            15'd31184: log10_cal = 16'b0000010111101111;
            15'd31185: log10_cal = 16'b0000010111101111;
            15'd31186: log10_cal = 16'b0000010111101111;
            15'd31187: log10_cal = 16'b0000010111101111;
            15'd31188: log10_cal = 16'b0000010111101111;
            15'd31189: log10_cal = 16'b0000010111101111;
            15'd31190: log10_cal = 16'b0000010111101111;
            15'd31191: log10_cal = 16'b0000010111101111;
            15'd31192: log10_cal = 16'b0000010111101111;
            15'd31193: log10_cal = 16'b0000010111101111;
            15'd31194: log10_cal = 16'b0000010111101111;
            15'd31195: log10_cal = 16'b0000010111101111;
            15'd31196: log10_cal = 16'b0000010111101111;
            15'd31197: log10_cal = 16'b0000010111101111;
            15'd31198: log10_cal = 16'b0000010111101111;
            15'd31199: log10_cal = 16'b0000010111101111;
            15'd31200: log10_cal = 16'b0000010111101111;
            15'd31201: log10_cal = 16'b0000010111101111;
            15'd31202: log10_cal = 16'b0000010111101111;
            15'd31203: log10_cal = 16'b0000010111101111;
            15'd31204: log10_cal = 16'b0000010111101111;
            15'd31205: log10_cal = 16'b0000010111101111;
            15'd31206: log10_cal = 16'b0000010111101111;
            15'd31207: log10_cal = 16'b0000010111101111;
            15'd31208: log10_cal = 16'b0000010111101111;
            15'd31209: log10_cal = 16'b0000010111101111;
            15'd31210: log10_cal = 16'b0000010111101111;
            15'd31211: log10_cal = 16'b0000010111101111;
            15'd31212: log10_cal = 16'b0000010111101111;
            15'd31213: log10_cal = 16'b0000010111101111;
            15'd31214: log10_cal = 16'b0000010111101111;
            15'd31215: log10_cal = 16'b0000010111101111;
            15'd31216: log10_cal = 16'b0000010111101111;
            15'd31217: log10_cal = 16'b0000010111101111;
            15'd31218: log10_cal = 16'b0000010111101111;
            15'd31219: log10_cal = 16'b0000010111101111;
            15'd31220: log10_cal = 16'b0000010111101111;
            15'd31221: log10_cal = 16'b0000010111101111;
            15'd31222: log10_cal = 16'b0000010111101111;
            15'd31223: log10_cal = 16'b0000010111101111;
            15'd31224: log10_cal = 16'b0000010111101111;
            15'd31225: log10_cal = 16'b0000010111101111;
            15'd31226: log10_cal = 16'b0000010111101111;
            15'd31227: log10_cal = 16'b0000010111101111;
            15'd31228: log10_cal = 16'b0000010111101111;
            15'd31229: log10_cal = 16'b0000010111101111;
            15'd31230: log10_cal = 16'b0000010111101111;
            15'd31231: log10_cal = 16'b0000010111101111;
            15'd31232: log10_cal = 16'b0000010111101111;
            15'd31233: log10_cal = 16'b0000010111101111;
            15'd31234: log10_cal = 16'b0000010111101111;
            15'd31235: log10_cal = 16'b0000010111101111;
            15'd31236: log10_cal = 16'b0000010111101111;
            15'd31237: log10_cal = 16'b0000010111101111;
            15'd31238: log10_cal = 16'b0000010111110000;
            15'd31239: log10_cal = 16'b0000010111110000;
            15'd31240: log10_cal = 16'b0000010111110000;
            15'd31241: log10_cal = 16'b0000010111110000;
            15'd31242: log10_cal = 16'b0000010111110000;
            15'd31243: log10_cal = 16'b0000010111110000;
            15'd31244: log10_cal = 16'b0000010111110000;
            15'd31245: log10_cal = 16'b0000010111110000;
            15'd31246: log10_cal = 16'b0000010111110000;
            15'd31247: log10_cal = 16'b0000010111110000;
            15'd31248: log10_cal = 16'b0000010111110000;
            15'd31249: log10_cal = 16'b0000010111110000;
            15'd31250: log10_cal = 16'b0000010111110000;
            15'd31251: log10_cal = 16'b0000010111110000;
            15'd31252: log10_cal = 16'b0000010111110000;
            15'd31253: log10_cal = 16'b0000010111110000;
            15'd31254: log10_cal = 16'b0000010111110000;
            15'd31255: log10_cal = 16'b0000010111110000;
            15'd31256: log10_cal = 16'b0000010111110000;
            15'd31257: log10_cal = 16'b0000010111110000;
            15'd31258: log10_cal = 16'b0000010111110000;
            15'd31259: log10_cal = 16'b0000010111110000;
            15'd31260: log10_cal = 16'b0000010111110000;
            15'd31261: log10_cal = 16'b0000010111110000;
            15'd31262: log10_cal = 16'b0000010111110000;
            15'd31263: log10_cal = 16'b0000010111110000;
            15'd31264: log10_cal = 16'b0000010111110000;
            15'd31265: log10_cal = 16'b0000010111110000;
            15'd31266: log10_cal = 16'b0000010111110000;
            15'd31267: log10_cal = 16'b0000010111110000;
            15'd31268: log10_cal = 16'b0000010111110000;
            15'd31269: log10_cal = 16'b0000010111110000;
            15'd31270: log10_cal = 16'b0000010111110000;
            15'd31271: log10_cal = 16'b0000010111110000;
            15'd31272: log10_cal = 16'b0000010111110000;
            15'd31273: log10_cal = 16'b0000010111110000;
            15'd31274: log10_cal = 16'b0000010111110000;
            15'd31275: log10_cal = 16'b0000010111110000;
            15'd31276: log10_cal = 16'b0000010111110000;
            15'd31277: log10_cal = 16'b0000010111110000;
            15'd31278: log10_cal = 16'b0000010111110000;
            15'd31279: log10_cal = 16'b0000010111110000;
            15'd31280: log10_cal = 16'b0000010111110000;
            15'd31281: log10_cal = 16'b0000010111110000;
            15'd31282: log10_cal = 16'b0000010111110000;
            15'd31283: log10_cal = 16'b0000010111110000;
            15'd31284: log10_cal = 16'b0000010111110000;
            15'd31285: log10_cal = 16'b0000010111110000;
            15'd31286: log10_cal = 16'b0000010111110000;
            15'd31287: log10_cal = 16'b0000010111110000;
            15'd31288: log10_cal = 16'b0000010111110000;
            15'd31289: log10_cal = 16'b0000010111110000;
            15'd31290: log10_cal = 16'b0000010111110000;
            15'd31291: log10_cal = 16'b0000010111110000;
            15'd31292: log10_cal = 16'b0000010111110000;
            15'd31293: log10_cal = 16'b0000010111110000;
            15'd31294: log10_cal = 16'b0000010111110000;
            15'd31295: log10_cal = 16'b0000010111110000;
            15'd31296: log10_cal = 16'b0000010111110000;
            15'd31297: log10_cal = 16'b0000010111110000;
            15'd31298: log10_cal = 16'b0000010111110000;
            15'd31299: log10_cal = 16'b0000010111110000;
            15'd31300: log10_cal = 16'b0000010111110000;
            15'd31301: log10_cal = 16'b0000010111110000;
            15'd31302: log10_cal = 16'b0000010111110000;
            15'd31303: log10_cal = 16'b0000010111110000;
            15'd31304: log10_cal = 16'b0000010111110000;
            15'd31305: log10_cal = 16'b0000010111110000;
            15'd31306: log10_cal = 16'b0000010111110000;
            15'd31307: log10_cal = 16'b0000010111110000;
            15'd31308: log10_cal = 16'b0000010111110001;
            15'd31309: log10_cal = 16'b0000010111110001;
            15'd31310: log10_cal = 16'b0000010111110001;
            15'd31311: log10_cal = 16'b0000010111110001;
            15'd31312: log10_cal = 16'b0000010111110001;
            15'd31313: log10_cal = 16'b0000010111110001;
            15'd31314: log10_cal = 16'b0000010111110001;
            15'd31315: log10_cal = 16'b0000010111110001;
            15'd31316: log10_cal = 16'b0000010111110001;
            15'd31317: log10_cal = 16'b0000010111110001;
            15'd31318: log10_cal = 16'b0000010111110001;
            15'd31319: log10_cal = 16'b0000010111110001;
            15'd31320: log10_cal = 16'b0000010111110001;
            15'd31321: log10_cal = 16'b0000010111110001;
            15'd31322: log10_cal = 16'b0000010111110001;
            15'd31323: log10_cal = 16'b0000010111110001;
            15'd31324: log10_cal = 16'b0000010111110001;
            15'd31325: log10_cal = 16'b0000010111110001;
            15'd31326: log10_cal = 16'b0000010111110001;
            15'd31327: log10_cal = 16'b0000010111110001;
            15'd31328: log10_cal = 16'b0000010111110001;
            15'd31329: log10_cal = 16'b0000010111110001;
            15'd31330: log10_cal = 16'b0000010111110001;
            15'd31331: log10_cal = 16'b0000010111110001;
            15'd31332: log10_cal = 16'b0000010111110001;
            15'd31333: log10_cal = 16'b0000010111110001;
            15'd31334: log10_cal = 16'b0000010111110001;
            15'd31335: log10_cal = 16'b0000010111110001;
            15'd31336: log10_cal = 16'b0000010111110001;
            15'd31337: log10_cal = 16'b0000010111110001;
            15'd31338: log10_cal = 16'b0000010111110001;
            15'd31339: log10_cal = 16'b0000010111110001;
            15'd31340: log10_cal = 16'b0000010111110001;
            15'd31341: log10_cal = 16'b0000010111110001;
            15'd31342: log10_cal = 16'b0000010111110001;
            15'd31343: log10_cal = 16'b0000010111110001;
            15'd31344: log10_cal = 16'b0000010111110001;
            15'd31345: log10_cal = 16'b0000010111110001;
            15'd31346: log10_cal = 16'b0000010111110001;
            15'd31347: log10_cal = 16'b0000010111110001;
            15'd31348: log10_cal = 16'b0000010111110001;
            15'd31349: log10_cal = 16'b0000010111110001;
            15'd31350: log10_cal = 16'b0000010111110001;
            15'd31351: log10_cal = 16'b0000010111110001;
            15'd31352: log10_cal = 16'b0000010111110001;
            15'd31353: log10_cal = 16'b0000010111110001;
            15'd31354: log10_cal = 16'b0000010111110001;
            15'd31355: log10_cal = 16'b0000010111110001;
            15'd31356: log10_cal = 16'b0000010111110001;
            15'd31357: log10_cal = 16'b0000010111110001;
            15'd31358: log10_cal = 16'b0000010111110001;
            15'd31359: log10_cal = 16'b0000010111110001;
            15'd31360: log10_cal = 16'b0000010111110001;
            15'd31361: log10_cal = 16'b0000010111110001;
            15'd31362: log10_cal = 16'b0000010111110001;
            15'd31363: log10_cal = 16'b0000010111110001;
            15'd31364: log10_cal = 16'b0000010111110001;
            15'd31365: log10_cal = 16'b0000010111110001;
            15'd31366: log10_cal = 16'b0000010111110001;
            15'd31367: log10_cal = 16'b0000010111110001;
            15'd31368: log10_cal = 16'b0000010111110001;
            15'd31369: log10_cal = 16'b0000010111110001;
            15'd31370: log10_cal = 16'b0000010111110001;
            15'd31371: log10_cal = 16'b0000010111110001;
            15'd31372: log10_cal = 16'b0000010111110001;
            15'd31373: log10_cal = 16'b0000010111110001;
            15'd31374: log10_cal = 16'b0000010111110001;
            15'd31375: log10_cal = 16'b0000010111110001;
            15'd31376: log10_cal = 16'b0000010111110001;
            15'd31377: log10_cal = 16'b0000010111110001;
            15'd31378: log10_cal = 16'b0000010111110001;
            15'd31379: log10_cal = 16'b0000010111110010;
            15'd31380: log10_cal = 16'b0000010111110010;
            15'd31381: log10_cal = 16'b0000010111110010;
            15'd31382: log10_cal = 16'b0000010111110010;
            15'd31383: log10_cal = 16'b0000010111110010;
            15'd31384: log10_cal = 16'b0000010111110010;
            15'd31385: log10_cal = 16'b0000010111110010;
            15'd31386: log10_cal = 16'b0000010111110010;
            15'd31387: log10_cal = 16'b0000010111110010;
            15'd31388: log10_cal = 16'b0000010111110010;
            15'd31389: log10_cal = 16'b0000010111110010;
            15'd31390: log10_cal = 16'b0000010111110010;
            15'd31391: log10_cal = 16'b0000010111110010;
            15'd31392: log10_cal = 16'b0000010111110010;
            15'd31393: log10_cal = 16'b0000010111110010;
            15'd31394: log10_cal = 16'b0000010111110010;
            15'd31395: log10_cal = 16'b0000010111110010;
            15'd31396: log10_cal = 16'b0000010111110010;
            15'd31397: log10_cal = 16'b0000010111110010;
            15'd31398: log10_cal = 16'b0000010111110010;
            15'd31399: log10_cal = 16'b0000010111110010;
            15'd31400: log10_cal = 16'b0000010111110010;
            15'd31401: log10_cal = 16'b0000010111110010;
            15'd31402: log10_cal = 16'b0000010111110010;
            15'd31403: log10_cal = 16'b0000010111110010;
            15'd31404: log10_cal = 16'b0000010111110010;
            15'd31405: log10_cal = 16'b0000010111110010;
            15'd31406: log10_cal = 16'b0000010111110010;
            15'd31407: log10_cal = 16'b0000010111110010;
            15'd31408: log10_cal = 16'b0000010111110010;
            15'd31409: log10_cal = 16'b0000010111110010;
            15'd31410: log10_cal = 16'b0000010111110010;
            15'd31411: log10_cal = 16'b0000010111110010;
            15'd31412: log10_cal = 16'b0000010111110010;
            15'd31413: log10_cal = 16'b0000010111110010;
            15'd31414: log10_cal = 16'b0000010111110010;
            15'd31415: log10_cal = 16'b0000010111110010;
            15'd31416: log10_cal = 16'b0000010111110010;
            15'd31417: log10_cal = 16'b0000010111110010;
            15'd31418: log10_cal = 16'b0000010111110010;
            15'd31419: log10_cal = 16'b0000010111110010;
            15'd31420: log10_cal = 16'b0000010111110010;
            15'd31421: log10_cal = 16'b0000010111110010;
            15'd31422: log10_cal = 16'b0000010111110010;
            15'd31423: log10_cal = 16'b0000010111110010;
            15'd31424: log10_cal = 16'b0000010111110010;
            15'd31425: log10_cal = 16'b0000010111110010;
            15'd31426: log10_cal = 16'b0000010111110010;
            15'd31427: log10_cal = 16'b0000010111110010;
            15'd31428: log10_cal = 16'b0000010111110010;
            15'd31429: log10_cal = 16'b0000010111110010;
            15'd31430: log10_cal = 16'b0000010111110010;
            15'd31431: log10_cal = 16'b0000010111110010;
            15'd31432: log10_cal = 16'b0000010111110010;
            15'd31433: log10_cal = 16'b0000010111110010;
            15'd31434: log10_cal = 16'b0000010111110010;
            15'd31435: log10_cal = 16'b0000010111110010;
            15'd31436: log10_cal = 16'b0000010111110010;
            15'd31437: log10_cal = 16'b0000010111110010;
            15'd31438: log10_cal = 16'b0000010111110010;
            15'd31439: log10_cal = 16'b0000010111110010;
            15'd31440: log10_cal = 16'b0000010111110010;
            15'd31441: log10_cal = 16'b0000010111110010;
            15'd31442: log10_cal = 16'b0000010111110010;
            15'd31443: log10_cal = 16'b0000010111110010;
            15'd31444: log10_cal = 16'b0000010111110010;
            15'd31445: log10_cal = 16'b0000010111110010;
            15'd31446: log10_cal = 16'b0000010111110010;
            15'd31447: log10_cal = 16'b0000010111110010;
            15'd31448: log10_cal = 16'b0000010111110010;
            15'd31449: log10_cal = 16'b0000010111110011;
            15'd31450: log10_cal = 16'b0000010111110011;
            15'd31451: log10_cal = 16'b0000010111110011;
            15'd31452: log10_cal = 16'b0000010111110011;
            15'd31453: log10_cal = 16'b0000010111110011;
            15'd31454: log10_cal = 16'b0000010111110011;
            15'd31455: log10_cal = 16'b0000010111110011;
            15'd31456: log10_cal = 16'b0000010111110011;
            15'd31457: log10_cal = 16'b0000010111110011;
            15'd31458: log10_cal = 16'b0000010111110011;
            15'd31459: log10_cal = 16'b0000010111110011;
            15'd31460: log10_cal = 16'b0000010111110011;
            15'd31461: log10_cal = 16'b0000010111110011;
            15'd31462: log10_cal = 16'b0000010111110011;
            15'd31463: log10_cal = 16'b0000010111110011;
            15'd31464: log10_cal = 16'b0000010111110011;
            15'd31465: log10_cal = 16'b0000010111110011;
            15'd31466: log10_cal = 16'b0000010111110011;
            15'd31467: log10_cal = 16'b0000010111110011;
            15'd31468: log10_cal = 16'b0000010111110011;
            15'd31469: log10_cal = 16'b0000010111110011;
            15'd31470: log10_cal = 16'b0000010111110011;
            15'd31471: log10_cal = 16'b0000010111110011;
            15'd31472: log10_cal = 16'b0000010111110011;
            15'd31473: log10_cal = 16'b0000010111110011;
            15'd31474: log10_cal = 16'b0000010111110011;
            15'd31475: log10_cal = 16'b0000010111110011;
            15'd31476: log10_cal = 16'b0000010111110011;
            15'd31477: log10_cal = 16'b0000010111110011;
            15'd31478: log10_cal = 16'b0000010111110011;
            15'd31479: log10_cal = 16'b0000010111110011;
            15'd31480: log10_cal = 16'b0000010111110011;
            15'd31481: log10_cal = 16'b0000010111110011;
            15'd31482: log10_cal = 16'b0000010111110011;
            15'd31483: log10_cal = 16'b0000010111110011;
            15'd31484: log10_cal = 16'b0000010111110011;
            15'd31485: log10_cal = 16'b0000010111110011;
            15'd31486: log10_cal = 16'b0000010111110011;
            15'd31487: log10_cal = 16'b0000010111110011;
            15'd31488: log10_cal = 16'b0000010111110011;
            15'd31489: log10_cal = 16'b0000010111110011;
            15'd31490: log10_cal = 16'b0000010111110011;
            15'd31491: log10_cal = 16'b0000010111110011;
            15'd31492: log10_cal = 16'b0000010111110011;
            15'd31493: log10_cal = 16'b0000010111110011;
            15'd31494: log10_cal = 16'b0000010111110011;
            15'd31495: log10_cal = 16'b0000010111110011;
            15'd31496: log10_cal = 16'b0000010111110011;
            15'd31497: log10_cal = 16'b0000010111110011;
            15'd31498: log10_cal = 16'b0000010111110011;
            15'd31499: log10_cal = 16'b0000010111110011;
            15'd31500: log10_cal = 16'b0000010111110011;
            15'd31501: log10_cal = 16'b0000010111110011;
            15'd31502: log10_cal = 16'b0000010111110011;
            15'd31503: log10_cal = 16'b0000010111110011;
            15'd31504: log10_cal = 16'b0000010111110011;
            15'd31505: log10_cal = 16'b0000010111110011;
            15'd31506: log10_cal = 16'b0000010111110011;
            15'd31507: log10_cal = 16'b0000010111110011;
            15'd31508: log10_cal = 16'b0000010111110011;
            15'd31509: log10_cal = 16'b0000010111110011;
            15'd31510: log10_cal = 16'b0000010111110011;
            15'd31511: log10_cal = 16'b0000010111110011;
            15'd31512: log10_cal = 16'b0000010111110011;
            15'd31513: log10_cal = 16'b0000010111110011;
            15'd31514: log10_cal = 16'b0000010111110011;
            15'd31515: log10_cal = 16'b0000010111110011;
            15'd31516: log10_cal = 16'b0000010111110011;
            15'd31517: log10_cal = 16'b0000010111110011;
            15'd31518: log10_cal = 16'b0000010111110011;
            15'd31519: log10_cal = 16'b0000010111110011;
            15'd31520: log10_cal = 16'b0000010111110100;
            15'd31521: log10_cal = 16'b0000010111110100;
            15'd31522: log10_cal = 16'b0000010111110100;
            15'd31523: log10_cal = 16'b0000010111110100;
            15'd31524: log10_cal = 16'b0000010111110100;
            15'd31525: log10_cal = 16'b0000010111110100;
            15'd31526: log10_cal = 16'b0000010111110100;
            15'd31527: log10_cal = 16'b0000010111110100;
            15'd31528: log10_cal = 16'b0000010111110100;
            15'd31529: log10_cal = 16'b0000010111110100;
            15'd31530: log10_cal = 16'b0000010111110100;
            15'd31531: log10_cal = 16'b0000010111110100;
            15'd31532: log10_cal = 16'b0000010111110100;
            15'd31533: log10_cal = 16'b0000010111110100;
            15'd31534: log10_cal = 16'b0000010111110100;
            15'd31535: log10_cal = 16'b0000010111110100;
            15'd31536: log10_cal = 16'b0000010111110100;
            15'd31537: log10_cal = 16'b0000010111110100;
            15'd31538: log10_cal = 16'b0000010111110100;
            15'd31539: log10_cal = 16'b0000010111110100;
            15'd31540: log10_cal = 16'b0000010111110100;
            15'd31541: log10_cal = 16'b0000010111110100;
            15'd31542: log10_cal = 16'b0000010111110100;
            15'd31543: log10_cal = 16'b0000010111110100;
            15'd31544: log10_cal = 16'b0000010111110100;
            15'd31545: log10_cal = 16'b0000010111110100;
            15'd31546: log10_cal = 16'b0000010111110100;
            15'd31547: log10_cal = 16'b0000010111110100;
            15'd31548: log10_cal = 16'b0000010111110100;
            15'd31549: log10_cal = 16'b0000010111110100;
            15'd31550: log10_cal = 16'b0000010111110100;
            15'd31551: log10_cal = 16'b0000010111110100;
            15'd31552: log10_cal = 16'b0000010111110100;
            15'd31553: log10_cal = 16'b0000010111110100;
            15'd31554: log10_cal = 16'b0000010111110100;
            15'd31555: log10_cal = 16'b0000010111110100;
            15'd31556: log10_cal = 16'b0000010111110100;
            15'd31557: log10_cal = 16'b0000010111110100;
            15'd31558: log10_cal = 16'b0000010111110100;
            15'd31559: log10_cal = 16'b0000010111110100;
            15'd31560: log10_cal = 16'b0000010111110100;
            15'd31561: log10_cal = 16'b0000010111110100;
            15'd31562: log10_cal = 16'b0000010111110100;
            15'd31563: log10_cal = 16'b0000010111110100;
            15'd31564: log10_cal = 16'b0000010111110100;
            15'd31565: log10_cal = 16'b0000010111110100;
            15'd31566: log10_cal = 16'b0000010111110100;
            15'd31567: log10_cal = 16'b0000010111110100;
            15'd31568: log10_cal = 16'b0000010111110100;
            15'd31569: log10_cal = 16'b0000010111110100;
            15'd31570: log10_cal = 16'b0000010111110100;
            15'd31571: log10_cal = 16'b0000010111110100;
            15'd31572: log10_cal = 16'b0000010111110100;
            15'd31573: log10_cal = 16'b0000010111110100;
            15'd31574: log10_cal = 16'b0000010111110100;
            15'd31575: log10_cal = 16'b0000010111110100;
            15'd31576: log10_cal = 16'b0000010111110100;
            15'd31577: log10_cal = 16'b0000010111110100;
            15'd31578: log10_cal = 16'b0000010111110100;
            15'd31579: log10_cal = 16'b0000010111110100;
            15'd31580: log10_cal = 16'b0000010111110100;
            15'd31581: log10_cal = 16'b0000010111110100;
            15'd31582: log10_cal = 16'b0000010111110100;
            15'd31583: log10_cal = 16'b0000010111110100;
            15'd31584: log10_cal = 16'b0000010111110100;
            15'd31585: log10_cal = 16'b0000010111110100;
            15'd31586: log10_cal = 16'b0000010111110100;
            15'd31587: log10_cal = 16'b0000010111110100;
            15'd31588: log10_cal = 16'b0000010111110100;
            15'd31589: log10_cal = 16'b0000010111110100;
            15'd31590: log10_cal = 16'b0000010111110100;
            15'd31591: log10_cal = 16'b0000010111110101;
            15'd31592: log10_cal = 16'b0000010111110101;
            15'd31593: log10_cal = 16'b0000010111110101;
            15'd31594: log10_cal = 16'b0000010111110101;
            15'd31595: log10_cal = 16'b0000010111110101;
            15'd31596: log10_cal = 16'b0000010111110101;
            15'd31597: log10_cal = 16'b0000010111110101;
            15'd31598: log10_cal = 16'b0000010111110101;
            15'd31599: log10_cal = 16'b0000010111110101;
            15'd31600: log10_cal = 16'b0000010111110101;
            15'd31601: log10_cal = 16'b0000010111110101;
            15'd31602: log10_cal = 16'b0000010111110101;
            15'd31603: log10_cal = 16'b0000010111110101;
            15'd31604: log10_cal = 16'b0000010111110101;
            15'd31605: log10_cal = 16'b0000010111110101;
            15'd31606: log10_cal = 16'b0000010111110101;
            15'd31607: log10_cal = 16'b0000010111110101;
            15'd31608: log10_cal = 16'b0000010111110101;
            15'd31609: log10_cal = 16'b0000010111110101;
            15'd31610: log10_cal = 16'b0000010111110101;
            15'd31611: log10_cal = 16'b0000010111110101;
            15'd31612: log10_cal = 16'b0000010111110101;
            15'd31613: log10_cal = 16'b0000010111110101;
            15'd31614: log10_cal = 16'b0000010111110101;
            15'd31615: log10_cal = 16'b0000010111110101;
            15'd31616: log10_cal = 16'b0000010111110101;
            15'd31617: log10_cal = 16'b0000010111110101;
            15'd31618: log10_cal = 16'b0000010111110101;
            15'd31619: log10_cal = 16'b0000010111110101;
            15'd31620: log10_cal = 16'b0000010111110101;
            15'd31621: log10_cal = 16'b0000010111110101;
            15'd31622: log10_cal = 16'b0000010111110101;
            15'd31623: log10_cal = 16'b0000010111110101;
            15'd31624: log10_cal = 16'b0000010111110101;
            15'd31625: log10_cal = 16'b0000010111110101;
            15'd31626: log10_cal = 16'b0000010111110101;
            15'd31627: log10_cal = 16'b0000010111110101;
            15'd31628: log10_cal = 16'b0000010111110101;
            15'd31629: log10_cal = 16'b0000010111110101;
            15'd31630: log10_cal = 16'b0000010111110101;
            15'd31631: log10_cal = 16'b0000010111110101;
            15'd31632: log10_cal = 16'b0000010111110101;
            15'd31633: log10_cal = 16'b0000010111110101;
            15'd31634: log10_cal = 16'b0000010111110101;
            15'd31635: log10_cal = 16'b0000010111110101;
            15'd31636: log10_cal = 16'b0000010111110101;
            15'd31637: log10_cal = 16'b0000010111110101;
            15'd31638: log10_cal = 16'b0000010111110101;
            15'd31639: log10_cal = 16'b0000010111110101;
            15'd31640: log10_cal = 16'b0000010111110101;
            15'd31641: log10_cal = 16'b0000010111110101;
            15'd31642: log10_cal = 16'b0000010111110101;
            15'd31643: log10_cal = 16'b0000010111110101;
            15'd31644: log10_cal = 16'b0000010111110101;
            15'd31645: log10_cal = 16'b0000010111110101;
            15'd31646: log10_cal = 16'b0000010111110101;
            15'd31647: log10_cal = 16'b0000010111110101;
            15'd31648: log10_cal = 16'b0000010111110101;
            15'd31649: log10_cal = 16'b0000010111110101;
            15'd31650: log10_cal = 16'b0000010111110101;
            15'd31651: log10_cal = 16'b0000010111110101;
            15'd31652: log10_cal = 16'b0000010111110101;
            15'd31653: log10_cal = 16'b0000010111110101;
            15'd31654: log10_cal = 16'b0000010111110101;
            15'd31655: log10_cal = 16'b0000010111110101;
            15'd31656: log10_cal = 16'b0000010111110101;
            15'd31657: log10_cal = 16'b0000010111110101;
            15'd31658: log10_cal = 16'b0000010111110101;
            15'd31659: log10_cal = 16'b0000010111110101;
            15'd31660: log10_cal = 16'b0000010111110101;
            15'd31661: log10_cal = 16'b0000010111110101;
            15'd31662: log10_cal = 16'b0000010111110110;
            15'd31663: log10_cal = 16'b0000010111110110;
            15'd31664: log10_cal = 16'b0000010111110110;
            15'd31665: log10_cal = 16'b0000010111110110;
            15'd31666: log10_cal = 16'b0000010111110110;
            15'd31667: log10_cal = 16'b0000010111110110;
            15'd31668: log10_cal = 16'b0000010111110110;
            15'd31669: log10_cal = 16'b0000010111110110;
            15'd31670: log10_cal = 16'b0000010111110110;
            15'd31671: log10_cal = 16'b0000010111110110;
            15'd31672: log10_cal = 16'b0000010111110110;
            15'd31673: log10_cal = 16'b0000010111110110;
            15'd31674: log10_cal = 16'b0000010111110110;
            15'd31675: log10_cal = 16'b0000010111110110;
            15'd31676: log10_cal = 16'b0000010111110110;
            15'd31677: log10_cal = 16'b0000010111110110;
            15'd31678: log10_cal = 16'b0000010111110110;
            15'd31679: log10_cal = 16'b0000010111110110;
            15'd31680: log10_cal = 16'b0000010111110110;
            15'd31681: log10_cal = 16'b0000010111110110;
            15'd31682: log10_cal = 16'b0000010111110110;
            15'd31683: log10_cal = 16'b0000010111110110;
            15'd31684: log10_cal = 16'b0000010111110110;
            15'd31685: log10_cal = 16'b0000010111110110;
            15'd31686: log10_cal = 16'b0000010111110110;
            15'd31687: log10_cal = 16'b0000010111110110;
            15'd31688: log10_cal = 16'b0000010111110110;
            15'd31689: log10_cal = 16'b0000010111110110;
            15'd31690: log10_cal = 16'b0000010111110110;
            15'd31691: log10_cal = 16'b0000010111110110;
            15'd31692: log10_cal = 16'b0000010111110110;
            15'd31693: log10_cal = 16'b0000010111110110;
            15'd31694: log10_cal = 16'b0000010111110110;
            15'd31695: log10_cal = 16'b0000010111110110;
            15'd31696: log10_cal = 16'b0000010111110110;
            15'd31697: log10_cal = 16'b0000010111110110;
            15'd31698: log10_cal = 16'b0000010111110110;
            15'd31699: log10_cal = 16'b0000010111110110;
            15'd31700: log10_cal = 16'b0000010111110110;
            15'd31701: log10_cal = 16'b0000010111110110;
            15'd31702: log10_cal = 16'b0000010111110110;
            15'd31703: log10_cal = 16'b0000010111110110;
            15'd31704: log10_cal = 16'b0000010111110110;
            15'd31705: log10_cal = 16'b0000010111110110;
            15'd31706: log10_cal = 16'b0000010111110110;
            15'd31707: log10_cal = 16'b0000010111110110;
            15'd31708: log10_cal = 16'b0000010111110110;
            15'd31709: log10_cal = 16'b0000010111110110;
            15'd31710: log10_cal = 16'b0000010111110110;
            15'd31711: log10_cal = 16'b0000010111110110;
            15'd31712: log10_cal = 16'b0000010111110110;
            15'd31713: log10_cal = 16'b0000010111110110;
            15'd31714: log10_cal = 16'b0000010111110110;
            15'd31715: log10_cal = 16'b0000010111110110;
            15'd31716: log10_cal = 16'b0000010111110110;
            15'd31717: log10_cal = 16'b0000010111110110;
            15'd31718: log10_cal = 16'b0000010111110110;
            15'd31719: log10_cal = 16'b0000010111110110;
            15'd31720: log10_cal = 16'b0000010111110110;
            15'd31721: log10_cal = 16'b0000010111110110;
            15'd31722: log10_cal = 16'b0000010111110110;
            15'd31723: log10_cal = 16'b0000010111110110;
            15'd31724: log10_cal = 16'b0000010111110110;
            15'd31725: log10_cal = 16'b0000010111110110;
            15'd31726: log10_cal = 16'b0000010111110110;
            15'd31727: log10_cal = 16'b0000010111110110;
            15'd31728: log10_cal = 16'b0000010111110110;
            15'd31729: log10_cal = 16'b0000010111110110;
            15'd31730: log10_cal = 16'b0000010111110110;
            15'd31731: log10_cal = 16'b0000010111110110;
            15'd31732: log10_cal = 16'b0000010111110110;
            15'd31733: log10_cal = 16'b0000010111110111;
            15'd31734: log10_cal = 16'b0000010111110111;
            15'd31735: log10_cal = 16'b0000010111110111;
            15'd31736: log10_cal = 16'b0000010111110111;
            15'd31737: log10_cal = 16'b0000010111110111;
            15'd31738: log10_cal = 16'b0000010111110111;
            15'd31739: log10_cal = 16'b0000010111110111;
            15'd31740: log10_cal = 16'b0000010111110111;
            15'd31741: log10_cal = 16'b0000010111110111;
            15'd31742: log10_cal = 16'b0000010111110111;
            15'd31743: log10_cal = 16'b0000010111110111;
            15'd31744: log10_cal = 16'b0000010111110111;
            15'd31745: log10_cal = 16'b0000010111110111;
            15'd31746: log10_cal = 16'b0000010111110111;
            15'd31747: log10_cal = 16'b0000010111110111;
            15'd31748: log10_cal = 16'b0000010111110111;
            15'd31749: log10_cal = 16'b0000010111110111;
            15'd31750: log10_cal = 16'b0000010111110111;
            15'd31751: log10_cal = 16'b0000010111110111;
            15'd31752: log10_cal = 16'b0000010111110111;
            15'd31753: log10_cal = 16'b0000010111110111;
            15'd31754: log10_cal = 16'b0000010111110111;
            15'd31755: log10_cal = 16'b0000010111110111;
            15'd31756: log10_cal = 16'b0000010111110111;
            15'd31757: log10_cal = 16'b0000010111110111;
            15'd31758: log10_cal = 16'b0000010111110111;
            15'd31759: log10_cal = 16'b0000010111110111;
            15'd31760: log10_cal = 16'b0000010111110111;
            15'd31761: log10_cal = 16'b0000010111110111;
            15'd31762: log10_cal = 16'b0000010111110111;
            15'd31763: log10_cal = 16'b0000010111110111;
            15'd31764: log10_cal = 16'b0000010111110111;
            15'd31765: log10_cal = 16'b0000010111110111;
            15'd31766: log10_cal = 16'b0000010111110111;
            15'd31767: log10_cal = 16'b0000010111110111;
            15'd31768: log10_cal = 16'b0000010111110111;
            15'd31769: log10_cal = 16'b0000010111110111;
            15'd31770: log10_cal = 16'b0000010111110111;
            15'd31771: log10_cal = 16'b0000010111110111;
            15'd31772: log10_cal = 16'b0000010111110111;
            15'd31773: log10_cal = 16'b0000010111110111;
            15'd31774: log10_cal = 16'b0000010111110111;
            15'd31775: log10_cal = 16'b0000010111110111;
            15'd31776: log10_cal = 16'b0000010111110111;
            15'd31777: log10_cal = 16'b0000010111110111;
            15'd31778: log10_cal = 16'b0000010111110111;
            15'd31779: log10_cal = 16'b0000010111110111;
            15'd31780: log10_cal = 16'b0000010111110111;
            15'd31781: log10_cal = 16'b0000010111110111;
            15'd31782: log10_cal = 16'b0000010111110111;
            15'd31783: log10_cal = 16'b0000010111110111;
            15'd31784: log10_cal = 16'b0000010111110111;
            15'd31785: log10_cal = 16'b0000010111110111;
            15'd31786: log10_cal = 16'b0000010111110111;
            15'd31787: log10_cal = 16'b0000010111110111;
            15'd31788: log10_cal = 16'b0000010111110111;
            15'd31789: log10_cal = 16'b0000010111110111;
            15'd31790: log10_cal = 16'b0000010111110111;
            15'd31791: log10_cal = 16'b0000010111110111;
            15'd31792: log10_cal = 16'b0000010111110111;
            15'd31793: log10_cal = 16'b0000010111110111;
            15'd31794: log10_cal = 16'b0000010111110111;
            15'd31795: log10_cal = 16'b0000010111110111;
            15'd31796: log10_cal = 16'b0000010111110111;
            15'd31797: log10_cal = 16'b0000010111110111;
            15'd31798: log10_cal = 16'b0000010111110111;
            15'd31799: log10_cal = 16'b0000010111110111;
            15'd31800: log10_cal = 16'b0000010111110111;
            15'd31801: log10_cal = 16'b0000010111110111;
            15'd31802: log10_cal = 16'b0000010111110111;
            15'd31803: log10_cal = 16'b0000010111110111;
            15'd31804: log10_cal = 16'b0000010111110111;
            15'd31805: log10_cal = 16'b0000010111111000;
            15'd31806: log10_cal = 16'b0000010111111000;
            15'd31807: log10_cal = 16'b0000010111111000;
            15'd31808: log10_cal = 16'b0000010111111000;
            15'd31809: log10_cal = 16'b0000010111111000;
            15'd31810: log10_cal = 16'b0000010111111000;
            15'd31811: log10_cal = 16'b0000010111111000;
            15'd31812: log10_cal = 16'b0000010111111000;
            15'd31813: log10_cal = 16'b0000010111111000;
            15'd31814: log10_cal = 16'b0000010111111000;
            15'd31815: log10_cal = 16'b0000010111111000;
            15'd31816: log10_cal = 16'b0000010111111000;
            15'd31817: log10_cal = 16'b0000010111111000;
            15'd31818: log10_cal = 16'b0000010111111000;
            15'd31819: log10_cal = 16'b0000010111111000;
            15'd31820: log10_cal = 16'b0000010111111000;
            15'd31821: log10_cal = 16'b0000010111111000;
            15'd31822: log10_cal = 16'b0000010111111000;
            15'd31823: log10_cal = 16'b0000010111111000;
            15'd31824: log10_cal = 16'b0000010111111000;
            15'd31825: log10_cal = 16'b0000010111111000;
            15'd31826: log10_cal = 16'b0000010111111000;
            15'd31827: log10_cal = 16'b0000010111111000;
            15'd31828: log10_cal = 16'b0000010111111000;
            15'd31829: log10_cal = 16'b0000010111111000;
            15'd31830: log10_cal = 16'b0000010111111000;
            15'd31831: log10_cal = 16'b0000010111111000;
            15'd31832: log10_cal = 16'b0000010111111000;
            15'd31833: log10_cal = 16'b0000010111111000;
            15'd31834: log10_cal = 16'b0000010111111000;
            15'd31835: log10_cal = 16'b0000010111111000;
            15'd31836: log10_cal = 16'b0000010111111000;
            15'd31837: log10_cal = 16'b0000010111111000;
            15'd31838: log10_cal = 16'b0000010111111000;
            15'd31839: log10_cal = 16'b0000010111111000;
            15'd31840: log10_cal = 16'b0000010111111000;
            15'd31841: log10_cal = 16'b0000010111111000;
            15'd31842: log10_cal = 16'b0000010111111000;
            15'd31843: log10_cal = 16'b0000010111111000;
            15'd31844: log10_cal = 16'b0000010111111000;
            15'd31845: log10_cal = 16'b0000010111111000;
            15'd31846: log10_cal = 16'b0000010111111000;
            15'd31847: log10_cal = 16'b0000010111111000;
            15'd31848: log10_cal = 16'b0000010111111000;
            15'd31849: log10_cal = 16'b0000010111111000;
            15'd31850: log10_cal = 16'b0000010111111000;
            15'd31851: log10_cal = 16'b0000010111111000;
            15'd31852: log10_cal = 16'b0000010111111000;
            15'd31853: log10_cal = 16'b0000010111111000;
            15'd31854: log10_cal = 16'b0000010111111000;
            15'd31855: log10_cal = 16'b0000010111111000;
            15'd31856: log10_cal = 16'b0000010111111000;
            15'd31857: log10_cal = 16'b0000010111111000;
            15'd31858: log10_cal = 16'b0000010111111000;
            15'd31859: log10_cal = 16'b0000010111111000;
            15'd31860: log10_cal = 16'b0000010111111000;
            15'd31861: log10_cal = 16'b0000010111111000;
            15'd31862: log10_cal = 16'b0000010111111000;
            15'd31863: log10_cal = 16'b0000010111111000;
            15'd31864: log10_cal = 16'b0000010111111000;
            15'd31865: log10_cal = 16'b0000010111111000;
            15'd31866: log10_cal = 16'b0000010111111000;
            15'd31867: log10_cal = 16'b0000010111111000;
            15'd31868: log10_cal = 16'b0000010111111000;
            15'd31869: log10_cal = 16'b0000010111111000;
            15'd31870: log10_cal = 16'b0000010111111000;
            15'd31871: log10_cal = 16'b0000010111111000;
            15'd31872: log10_cal = 16'b0000010111111000;
            15'd31873: log10_cal = 16'b0000010111111000;
            15'd31874: log10_cal = 16'b0000010111111000;
            15'd31875: log10_cal = 16'b0000010111111000;
            15'd31876: log10_cal = 16'b0000010111111000;
            15'd31877: log10_cal = 16'b0000010111111001;
            15'd31878: log10_cal = 16'b0000010111111001;
            15'd31879: log10_cal = 16'b0000010111111001;
            15'd31880: log10_cal = 16'b0000010111111001;
            15'd31881: log10_cal = 16'b0000010111111001;
            15'd31882: log10_cal = 16'b0000010111111001;
            15'd31883: log10_cal = 16'b0000010111111001;
            15'd31884: log10_cal = 16'b0000010111111001;
            15'd31885: log10_cal = 16'b0000010111111001;
            15'd31886: log10_cal = 16'b0000010111111001;
            15'd31887: log10_cal = 16'b0000010111111001;
            15'd31888: log10_cal = 16'b0000010111111001;
            15'd31889: log10_cal = 16'b0000010111111001;
            15'd31890: log10_cal = 16'b0000010111111001;
            15'd31891: log10_cal = 16'b0000010111111001;
            15'd31892: log10_cal = 16'b0000010111111001;
            15'd31893: log10_cal = 16'b0000010111111001;
            15'd31894: log10_cal = 16'b0000010111111001;
            15'd31895: log10_cal = 16'b0000010111111001;
            15'd31896: log10_cal = 16'b0000010111111001;
            15'd31897: log10_cal = 16'b0000010111111001;
            15'd31898: log10_cal = 16'b0000010111111001;
            15'd31899: log10_cal = 16'b0000010111111001;
            15'd31900: log10_cal = 16'b0000010111111001;
            15'd31901: log10_cal = 16'b0000010111111001;
            15'd31902: log10_cal = 16'b0000010111111001;
            15'd31903: log10_cal = 16'b0000010111111001;
            15'd31904: log10_cal = 16'b0000010111111001;
            15'd31905: log10_cal = 16'b0000010111111001;
            15'd31906: log10_cal = 16'b0000010111111001;
            15'd31907: log10_cal = 16'b0000010111111001;
            15'd31908: log10_cal = 16'b0000010111111001;
            15'd31909: log10_cal = 16'b0000010111111001;
            15'd31910: log10_cal = 16'b0000010111111001;
            15'd31911: log10_cal = 16'b0000010111111001;
            15'd31912: log10_cal = 16'b0000010111111001;
            15'd31913: log10_cal = 16'b0000010111111001;
            15'd31914: log10_cal = 16'b0000010111111001;
            15'd31915: log10_cal = 16'b0000010111111001;
            15'd31916: log10_cal = 16'b0000010111111001;
            15'd31917: log10_cal = 16'b0000010111111001;
            15'd31918: log10_cal = 16'b0000010111111001;
            15'd31919: log10_cal = 16'b0000010111111001;
            15'd31920: log10_cal = 16'b0000010111111001;
            15'd31921: log10_cal = 16'b0000010111111001;
            15'd31922: log10_cal = 16'b0000010111111001;
            15'd31923: log10_cal = 16'b0000010111111001;
            15'd31924: log10_cal = 16'b0000010111111001;
            15'd31925: log10_cal = 16'b0000010111111001;
            15'd31926: log10_cal = 16'b0000010111111001;
            15'd31927: log10_cal = 16'b0000010111111001;
            15'd31928: log10_cal = 16'b0000010111111001;
            15'd31929: log10_cal = 16'b0000010111111001;
            15'd31930: log10_cal = 16'b0000010111111001;
            15'd31931: log10_cal = 16'b0000010111111001;
            15'd31932: log10_cal = 16'b0000010111111001;
            15'd31933: log10_cal = 16'b0000010111111001;
            15'd31934: log10_cal = 16'b0000010111111001;
            15'd31935: log10_cal = 16'b0000010111111001;
            15'd31936: log10_cal = 16'b0000010111111001;
            15'd31937: log10_cal = 16'b0000010111111001;
            15'd31938: log10_cal = 16'b0000010111111001;
            15'd31939: log10_cal = 16'b0000010111111001;
            15'd31940: log10_cal = 16'b0000010111111001;
            15'd31941: log10_cal = 16'b0000010111111001;
            15'd31942: log10_cal = 16'b0000010111111001;
            15'd31943: log10_cal = 16'b0000010111111001;
            15'd31944: log10_cal = 16'b0000010111111001;
            15'd31945: log10_cal = 16'b0000010111111001;
            15'd31946: log10_cal = 16'b0000010111111001;
            15'd31947: log10_cal = 16'b0000010111111001;
            15'd31948: log10_cal = 16'b0000010111111010;
            15'd31949: log10_cal = 16'b0000010111111010;
            15'd31950: log10_cal = 16'b0000010111111010;
            15'd31951: log10_cal = 16'b0000010111111010;
            15'd31952: log10_cal = 16'b0000010111111010;
            15'd31953: log10_cal = 16'b0000010111111010;
            15'd31954: log10_cal = 16'b0000010111111010;
            15'd31955: log10_cal = 16'b0000010111111010;
            15'd31956: log10_cal = 16'b0000010111111010;
            15'd31957: log10_cal = 16'b0000010111111010;
            15'd31958: log10_cal = 16'b0000010111111010;
            15'd31959: log10_cal = 16'b0000010111111010;
            15'd31960: log10_cal = 16'b0000010111111010;
            15'd31961: log10_cal = 16'b0000010111111010;
            15'd31962: log10_cal = 16'b0000010111111010;
            15'd31963: log10_cal = 16'b0000010111111010;
            15'd31964: log10_cal = 16'b0000010111111010;
            15'd31965: log10_cal = 16'b0000010111111010;
            15'd31966: log10_cal = 16'b0000010111111010;
            15'd31967: log10_cal = 16'b0000010111111010;
            15'd31968: log10_cal = 16'b0000010111111010;
            15'd31969: log10_cal = 16'b0000010111111010;
            15'd31970: log10_cal = 16'b0000010111111010;
            15'd31971: log10_cal = 16'b0000010111111010;
            15'd31972: log10_cal = 16'b0000010111111010;
            15'd31973: log10_cal = 16'b0000010111111010;
            15'd31974: log10_cal = 16'b0000010111111010;
            15'd31975: log10_cal = 16'b0000010111111010;
            15'd31976: log10_cal = 16'b0000010111111010;
            15'd31977: log10_cal = 16'b0000010111111010;
            15'd31978: log10_cal = 16'b0000010111111010;
            15'd31979: log10_cal = 16'b0000010111111010;
            15'd31980: log10_cal = 16'b0000010111111010;
            15'd31981: log10_cal = 16'b0000010111111010;
            15'd31982: log10_cal = 16'b0000010111111010;
            15'd31983: log10_cal = 16'b0000010111111010;
            15'd31984: log10_cal = 16'b0000010111111010;
            15'd31985: log10_cal = 16'b0000010111111010;
            15'd31986: log10_cal = 16'b0000010111111010;
            15'd31987: log10_cal = 16'b0000010111111010;
            15'd31988: log10_cal = 16'b0000010111111010;
            15'd31989: log10_cal = 16'b0000010111111010;
            15'd31990: log10_cal = 16'b0000010111111010;
            15'd31991: log10_cal = 16'b0000010111111010;
            15'd31992: log10_cal = 16'b0000010111111010;
            15'd31993: log10_cal = 16'b0000010111111010;
            15'd31994: log10_cal = 16'b0000010111111010;
            15'd31995: log10_cal = 16'b0000010111111010;
            15'd31996: log10_cal = 16'b0000010111111010;
            15'd31997: log10_cal = 16'b0000010111111010;
            15'd31998: log10_cal = 16'b0000010111111010;
            15'd31999: log10_cal = 16'b0000010111111010;
            15'd32000: log10_cal = 16'b0000010111111010;
            15'd32001: log10_cal = 16'b0000010111111010;
            15'd32002: log10_cal = 16'b0000010111111010;
            15'd32003: log10_cal = 16'b0000010111111010;
            15'd32004: log10_cal = 16'b0000010111111010;
            15'd32005: log10_cal = 16'b0000010111111010;
            15'd32006: log10_cal = 16'b0000010111111010;
            15'd32007: log10_cal = 16'b0000010111111010;
            15'd32008: log10_cal = 16'b0000010111111010;
            15'd32009: log10_cal = 16'b0000010111111010;
            15'd32010: log10_cal = 16'b0000010111111010;
            15'd32011: log10_cal = 16'b0000010111111010;
            15'd32012: log10_cal = 16'b0000010111111010;
            15'd32013: log10_cal = 16'b0000010111111010;
            15'd32014: log10_cal = 16'b0000010111111010;
            15'd32015: log10_cal = 16'b0000010111111010;
            15'd32016: log10_cal = 16'b0000010111111010;
            15'd32017: log10_cal = 16'b0000010111111010;
            15'd32018: log10_cal = 16'b0000010111111010;
            15'd32019: log10_cal = 16'b0000010111111010;
            15'd32020: log10_cal = 16'b0000010111111011;
            15'd32021: log10_cal = 16'b0000010111111011;
            15'd32022: log10_cal = 16'b0000010111111011;
            15'd32023: log10_cal = 16'b0000010111111011;
            15'd32024: log10_cal = 16'b0000010111111011;
            15'd32025: log10_cal = 16'b0000010111111011;
            15'd32026: log10_cal = 16'b0000010111111011;
            15'd32027: log10_cal = 16'b0000010111111011;
            15'd32028: log10_cal = 16'b0000010111111011;
            15'd32029: log10_cal = 16'b0000010111111011;
            15'd32030: log10_cal = 16'b0000010111111011;
            15'd32031: log10_cal = 16'b0000010111111011;
            15'd32032: log10_cal = 16'b0000010111111011;
            15'd32033: log10_cal = 16'b0000010111111011;
            15'd32034: log10_cal = 16'b0000010111111011;
            15'd32035: log10_cal = 16'b0000010111111011;
            15'd32036: log10_cal = 16'b0000010111111011;
            15'd32037: log10_cal = 16'b0000010111111011;
            15'd32038: log10_cal = 16'b0000010111111011;
            15'd32039: log10_cal = 16'b0000010111111011;
            15'd32040: log10_cal = 16'b0000010111111011;
            15'd32041: log10_cal = 16'b0000010111111011;
            15'd32042: log10_cal = 16'b0000010111111011;
            15'd32043: log10_cal = 16'b0000010111111011;
            15'd32044: log10_cal = 16'b0000010111111011;
            15'd32045: log10_cal = 16'b0000010111111011;
            15'd32046: log10_cal = 16'b0000010111111011;
            15'd32047: log10_cal = 16'b0000010111111011;
            15'd32048: log10_cal = 16'b0000010111111011;
            15'd32049: log10_cal = 16'b0000010111111011;
            15'd32050: log10_cal = 16'b0000010111111011;
            15'd32051: log10_cal = 16'b0000010111111011;
            15'd32052: log10_cal = 16'b0000010111111011;
            15'd32053: log10_cal = 16'b0000010111111011;
            15'd32054: log10_cal = 16'b0000010111111011;
            15'd32055: log10_cal = 16'b0000010111111011;
            15'd32056: log10_cal = 16'b0000010111111011;
            15'd32057: log10_cal = 16'b0000010111111011;
            15'd32058: log10_cal = 16'b0000010111111011;
            15'd32059: log10_cal = 16'b0000010111111011;
            15'd32060: log10_cal = 16'b0000010111111011;
            15'd32061: log10_cal = 16'b0000010111111011;
            15'd32062: log10_cal = 16'b0000010111111011;
            15'd32063: log10_cal = 16'b0000010111111011;
            15'd32064: log10_cal = 16'b0000010111111011;
            15'd32065: log10_cal = 16'b0000010111111011;
            15'd32066: log10_cal = 16'b0000010111111011;
            15'd32067: log10_cal = 16'b0000010111111011;
            15'd32068: log10_cal = 16'b0000010111111011;
            15'd32069: log10_cal = 16'b0000010111111011;
            15'd32070: log10_cal = 16'b0000010111111011;
            15'd32071: log10_cal = 16'b0000010111111011;
            15'd32072: log10_cal = 16'b0000010111111011;
            15'd32073: log10_cal = 16'b0000010111111011;
            15'd32074: log10_cal = 16'b0000010111111011;
            15'd32075: log10_cal = 16'b0000010111111011;
            15'd32076: log10_cal = 16'b0000010111111011;
            15'd32077: log10_cal = 16'b0000010111111011;
            15'd32078: log10_cal = 16'b0000010111111011;
            15'd32079: log10_cal = 16'b0000010111111011;
            15'd32080: log10_cal = 16'b0000010111111011;
            15'd32081: log10_cal = 16'b0000010111111011;
            15'd32082: log10_cal = 16'b0000010111111011;
            15'd32083: log10_cal = 16'b0000010111111011;
            15'd32084: log10_cal = 16'b0000010111111011;
            15'd32085: log10_cal = 16'b0000010111111011;
            15'd32086: log10_cal = 16'b0000010111111011;
            15'd32087: log10_cal = 16'b0000010111111011;
            15'd32088: log10_cal = 16'b0000010111111011;
            15'd32089: log10_cal = 16'b0000010111111011;
            15'd32090: log10_cal = 16'b0000010111111011;
            15'd32091: log10_cal = 16'b0000010111111011;
            15'd32092: log10_cal = 16'b0000010111111100;
            15'd32093: log10_cal = 16'b0000010111111100;
            15'd32094: log10_cal = 16'b0000010111111100;
            15'd32095: log10_cal = 16'b0000010111111100;
            15'd32096: log10_cal = 16'b0000010111111100;
            15'd32097: log10_cal = 16'b0000010111111100;
            15'd32098: log10_cal = 16'b0000010111111100;
            15'd32099: log10_cal = 16'b0000010111111100;
            15'd32100: log10_cal = 16'b0000010111111100;
            15'd32101: log10_cal = 16'b0000010111111100;
            15'd32102: log10_cal = 16'b0000010111111100;
            15'd32103: log10_cal = 16'b0000010111111100;
            15'd32104: log10_cal = 16'b0000010111111100;
            15'd32105: log10_cal = 16'b0000010111111100;
            15'd32106: log10_cal = 16'b0000010111111100;
            15'd32107: log10_cal = 16'b0000010111111100;
            15'd32108: log10_cal = 16'b0000010111111100;
            15'd32109: log10_cal = 16'b0000010111111100;
            15'd32110: log10_cal = 16'b0000010111111100;
            15'd32111: log10_cal = 16'b0000010111111100;
            15'd32112: log10_cal = 16'b0000010111111100;
            15'd32113: log10_cal = 16'b0000010111111100;
            15'd32114: log10_cal = 16'b0000010111111100;
            15'd32115: log10_cal = 16'b0000010111111100;
            15'd32116: log10_cal = 16'b0000010111111100;
            15'd32117: log10_cal = 16'b0000010111111100;
            15'd32118: log10_cal = 16'b0000010111111100;
            15'd32119: log10_cal = 16'b0000010111111100;
            15'd32120: log10_cal = 16'b0000010111111100;
            15'd32121: log10_cal = 16'b0000010111111100;
            15'd32122: log10_cal = 16'b0000010111111100;
            15'd32123: log10_cal = 16'b0000010111111100;
            15'd32124: log10_cal = 16'b0000010111111100;
            15'd32125: log10_cal = 16'b0000010111111100;
            15'd32126: log10_cal = 16'b0000010111111100;
            15'd32127: log10_cal = 16'b0000010111111100;
            15'd32128: log10_cal = 16'b0000010111111100;
            15'd32129: log10_cal = 16'b0000010111111100;
            15'd32130: log10_cal = 16'b0000010111111100;
            15'd32131: log10_cal = 16'b0000010111111100;
            15'd32132: log10_cal = 16'b0000010111111100;
            15'd32133: log10_cal = 16'b0000010111111100;
            15'd32134: log10_cal = 16'b0000010111111100;
            15'd32135: log10_cal = 16'b0000010111111100;
            15'd32136: log10_cal = 16'b0000010111111100;
            15'd32137: log10_cal = 16'b0000010111111100;
            15'd32138: log10_cal = 16'b0000010111111100;
            15'd32139: log10_cal = 16'b0000010111111100;
            15'd32140: log10_cal = 16'b0000010111111100;
            15'd32141: log10_cal = 16'b0000010111111100;
            15'd32142: log10_cal = 16'b0000010111111100;
            15'd32143: log10_cal = 16'b0000010111111100;
            15'd32144: log10_cal = 16'b0000010111111100;
            15'd32145: log10_cal = 16'b0000010111111100;
            15'd32146: log10_cal = 16'b0000010111111100;
            15'd32147: log10_cal = 16'b0000010111111100;
            15'd32148: log10_cal = 16'b0000010111111100;
            15'd32149: log10_cal = 16'b0000010111111100;
            15'd32150: log10_cal = 16'b0000010111111100;
            15'd32151: log10_cal = 16'b0000010111111100;
            15'd32152: log10_cal = 16'b0000010111111100;
            15'd32153: log10_cal = 16'b0000010111111100;
            15'd32154: log10_cal = 16'b0000010111111100;
            15'd32155: log10_cal = 16'b0000010111111100;
            15'd32156: log10_cal = 16'b0000010111111100;
            15'd32157: log10_cal = 16'b0000010111111100;
            15'd32158: log10_cal = 16'b0000010111111100;
            15'd32159: log10_cal = 16'b0000010111111100;
            15'd32160: log10_cal = 16'b0000010111111100;
            15'd32161: log10_cal = 16'b0000010111111100;
            15'd32162: log10_cal = 16'b0000010111111100;
            15'd32163: log10_cal = 16'b0000010111111100;
            15'd32164: log10_cal = 16'b0000010111111100;
            15'd32165: log10_cal = 16'b0000010111111101;
            15'd32166: log10_cal = 16'b0000010111111101;
            15'd32167: log10_cal = 16'b0000010111111101;
            15'd32168: log10_cal = 16'b0000010111111101;
            15'd32169: log10_cal = 16'b0000010111111101;
            15'd32170: log10_cal = 16'b0000010111111101;
            15'd32171: log10_cal = 16'b0000010111111101;
            15'd32172: log10_cal = 16'b0000010111111101;
            15'd32173: log10_cal = 16'b0000010111111101;
            15'd32174: log10_cal = 16'b0000010111111101;
            15'd32175: log10_cal = 16'b0000010111111101;
            15'd32176: log10_cal = 16'b0000010111111101;
            15'd32177: log10_cal = 16'b0000010111111101;
            15'd32178: log10_cal = 16'b0000010111111101;
            15'd32179: log10_cal = 16'b0000010111111101;
            15'd32180: log10_cal = 16'b0000010111111101;
            15'd32181: log10_cal = 16'b0000010111111101;
            15'd32182: log10_cal = 16'b0000010111111101;
            15'd32183: log10_cal = 16'b0000010111111101;
            15'd32184: log10_cal = 16'b0000010111111101;
            15'd32185: log10_cal = 16'b0000010111111101;
            15'd32186: log10_cal = 16'b0000010111111101;
            15'd32187: log10_cal = 16'b0000010111111101;
            15'd32188: log10_cal = 16'b0000010111111101;
            15'd32189: log10_cal = 16'b0000010111111101;
            15'd32190: log10_cal = 16'b0000010111111101;
            15'd32191: log10_cal = 16'b0000010111111101;
            15'd32192: log10_cal = 16'b0000010111111101;
            15'd32193: log10_cal = 16'b0000010111111101;
            15'd32194: log10_cal = 16'b0000010111111101;
            15'd32195: log10_cal = 16'b0000010111111101;
            15'd32196: log10_cal = 16'b0000010111111101;
            15'd32197: log10_cal = 16'b0000010111111101;
            15'd32198: log10_cal = 16'b0000010111111101;
            15'd32199: log10_cal = 16'b0000010111111101;
            15'd32200: log10_cal = 16'b0000010111111101;
            15'd32201: log10_cal = 16'b0000010111111101;
            15'd32202: log10_cal = 16'b0000010111111101;
            15'd32203: log10_cal = 16'b0000010111111101;
            15'd32204: log10_cal = 16'b0000010111111101;
            15'd32205: log10_cal = 16'b0000010111111101;
            15'd32206: log10_cal = 16'b0000010111111101;
            15'd32207: log10_cal = 16'b0000010111111101;
            15'd32208: log10_cal = 16'b0000010111111101;
            15'd32209: log10_cal = 16'b0000010111111101;
            15'd32210: log10_cal = 16'b0000010111111101;
            15'd32211: log10_cal = 16'b0000010111111101;
            15'd32212: log10_cal = 16'b0000010111111101;
            15'd32213: log10_cal = 16'b0000010111111101;
            15'd32214: log10_cal = 16'b0000010111111101;
            15'd32215: log10_cal = 16'b0000010111111101;
            15'd32216: log10_cal = 16'b0000010111111101;
            15'd32217: log10_cal = 16'b0000010111111101;
            15'd32218: log10_cal = 16'b0000010111111101;
            15'd32219: log10_cal = 16'b0000010111111101;
            15'd32220: log10_cal = 16'b0000010111111101;
            15'd32221: log10_cal = 16'b0000010111111101;
            15'd32222: log10_cal = 16'b0000010111111101;
            15'd32223: log10_cal = 16'b0000010111111101;
            15'd32224: log10_cal = 16'b0000010111111101;
            15'd32225: log10_cal = 16'b0000010111111101;
            15'd32226: log10_cal = 16'b0000010111111101;
            15'd32227: log10_cal = 16'b0000010111111101;
            15'd32228: log10_cal = 16'b0000010111111101;
            15'd32229: log10_cal = 16'b0000010111111101;
            15'd32230: log10_cal = 16'b0000010111111101;
            15'd32231: log10_cal = 16'b0000010111111101;
            15'd32232: log10_cal = 16'b0000010111111101;
            15'd32233: log10_cal = 16'b0000010111111101;
            15'd32234: log10_cal = 16'b0000010111111101;
            15'd32235: log10_cal = 16'b0000010111111101;
            15'd32236: log10_cal = 16'b0000010111111101;
            15'd32237: log10_cal = 16'b0000010111111110;
            15'd32238: log10_cal = 16'b0000010111111110;
            15'd32239: log10_cal = 16'b0000010111111110;
            15'd32240: log10_cal = 16'b0000010111111110;
            15'd32241: log10_cal = 16'b0000010111111110;
            15'd32242: log10_cal = 16'b0000010111111110;
            15'd32243: log10_cal = 16'b0000010111111110;
            15'd32244: log10_cal = 16'b0000010111111110;
            15'd32245: log10_cal = 16'b0000010111111110;
            15'd32246: log10_cal = 16'b0000010111111110;
            15'd32247: log10_cal = 16'b0000010111111110;
            15'd32248: log10_cal = 16'b0000010111111110;
            15'd32249: log10_cal = 16'b0000010111111110;
            15'd32250: log10_cal = 16'b0000010111111110;
            15'd32251: log10_cal = 16'b0000010111111110;
            15'd32252: log10_cal = 16'b0000010111111110;
            15'd32253: log10_cal = 16'b0000010111111110;
            15'd32254: log10_cal = 16'b0000010111111110;
            15'd32255: log10_cal = 16'b0000010111111110;
            15'd32256: log10_cal = 16'b0000010111111110;
            15'd32257: log10_cal = 16'b0000010111111110;
            15'd32258: log10_cal = 16'b0000010111111110;
            15'd32259: log10_cal = 16'b0000010111111110;
            15'd32260: log10_cal = 16'b0000010111111110;
            15'd32261: log10_cal = 16'b0000010111111110;
            15'd32262: log10_cal = 16'b0000010111111110;
            15'd32263: log10_cal = 16'b0000010111111110;
            15'd32264: log10_cal = 16'b0000010111111110;
            15'd32265: log10_cal = 16'b0000010111111110;
            15'd32266: log10_cal = 16'b0000010111111110;
            15'd32267: log10_cal = 16'b0000010111111110;
            15'd32268: log10_cal = 16'b0000010111111110;
            15'd32269: log10_cal = 16'b0000010111111110;
            15'd32270: log10_cal = 16'b0000010111111110;
            15'd32271: log10_cal = 16'b0000010111111110;
            15'd32272: log10_cal = 16'b0000010111111110;
            15'd32273: log10_cal = 16'b0000010111111110;
            15'd32274: log10_cal = 16'b0000010111111110;
            15'd32275: log10_cal = 16'b0000010111111110;
            15'd32276: log10_cal = 16'b0000010111111110;
            15'd32277: log10_cal = 16'b0000010111111110;
            15'd32278: log10_cal = 16'b0000010111111110;
            15'd32279: log10_cal = 16'b0000010111111110;
            15'd32280: log10_cal = 16'b0000010111111110;
            15'd32281: log10_cal = 16'b0000010111111110;
            15'd32282: log10_cal = 16'b0000010111111110;
            15'd32283: log10_cal = 16'b0000010111111110;
            15'd32284: log10_cal = 16'b0000010111111110;
            15'd32285: log10_cal = 16'b0000010111111110;
            15'd32286: log10_cal = 16'b0000010111111110;
            15'd32287: log10_cal = 16'b0000010111111110;
            15'd32288: log10_cal = 16'b0000010111111110;
            15'd32289: log10_cal = 16'b0000010111111110;
            15'd32290: log10_cal = 16'b0000010111111110;
            15'd32291: log10_cal = 16'b0000010111111110;
            15'd32292: log10_cal = 16'b0000010111111110;
            15'd32293: log10_cal = 16'b0000010111111110;
            15'd32294: log10_cal = 16'b0000010111111110;
            15'd32295: log10_cal = 16'b0000010111111110;
            15'd32296: log10_cal = 16'b0000010111111110;
            15'd32297: log10_cal = 16'b0000010111111110;
            15'd32298: log10_cal = 16'b0000010111111110;
            15'd32299: log10_cal = 16'b0000010111111110;
            15'd32300: log10_cal = 16'b0000010111111110;
            15'd32301: log10_cal = 16'b0000010111111110;
            15'd32302: log10_cal = 16'b0000010111111110;
            15'd32303: log10_cal = 16'b0000010111111110;
            15'd32304: log10_cal = 16'b0000010111111110;
            15'd32305: log10_cal = 16'b0000010111111110;
            15'd32306: log10_cal = 16'b0000010111111110;
            15'd32307: log10_cal = 16'b0000010111111110;
            15'd32308: log10_cal = 16'b0000010111111110;
            15'd32309: log10_cal = 16'b0000010111111111;
            15'd32310: log10_cal = 16'b0000010111111111;
            15'd32311: log10_cal = 16'b0000010111111111;
            15'd32312: log10_cal = 16'b0000010111111111;
            15'd32313: log10_cal = 16'b0000010111111111;
            15'd32314: log10_cal = 16'b0000010111111111;
            15'd32315: log10_cal = 16'b0000010111111111;
            15'd32316: log10_cal = 16'b0000010111111111;
            15'd32317: log10_cal = 16'b0000010111111111;
            15'd32318: log10_cal = 16'b0000010111111111;
            15'd32319: log10_cal = 16'b0000010111111111;
            15'd32320: log10_cal = 16'b0000010111111111;
            15'd32321: log10_cal = 16'b0000010111111111;
            15'd32322: log10_cal = 16'b0000010111111111;
            15'd32323: log10_cal = 16'b0000010111111111;
            15'd32324: log10_cal = 16'b0000010111111111;
            15'd32325: log10_cal = 16'b0000010111111111;
            15'd32326: log10_cal = 16'b0000010111111111;
            15'd32327: log10_cal = 16'b0000010111111111;
            15'd32328: log10_cal = 16'b0000010111111111;
            15'd32329: log10_cal = 16'b0000010111111111;
            15'd32330: log10_cal = 16'b0000010111111111;
            15'd32331: log10_cal = 16'b0000010111111111;
            15'd32332: log10_cal = 16'b0000010111111111;
            15'd32333: log10_cal = 16'b0000010111111111;
            15'd32334: log10_cal = 16'b0000010111111111;
            15'd32335: log10_cal = 16'b0000010111111111;
            15'd32336: log10_cal = 16'b0000010111111111;
            15'd32337: log10_cal = 16'b0000010111111111;
            15'd32338: log10_cal = 16'b0000010111111111;
            15'd32339: log10_cal = 16'b0000010111111111;
            15'd32340: log10_cal = 16'b0000010111111111;
            15'd32341: log10_cal = 16'b0000010111111111;
            15'd32342: log10_cal = 16'b0000010111111111;
            15'd32343: log10_cal = 16'b0000010111111111;
            15'd32344: log10_cal = 16'b0000010111111111;
            15'd32345: log10_cal = 16'b0000010111111111;
            15'd32346: log10_cal = 16'b0000010111111111;
            15'd32347: log10_cal = 16'b0000010111111111;
            15'd32348: log10_cal = 16'b0000010111111111;
            15'd32349: log10_cal = 16'b0000010111111111;
            15'd32350: log10_cal = 16'b0000010111111111;
            15'd32351: log10_cal = 16'b0000010111111111;
            15'd32352: log10_cal = 16'b0000010111111111;
            15'd32353: log10_cal = 16'b0000010111111111;
            15'd32354: log10_cal = 16'b0000010111111111;
            15'd32355: log10_cal = 16'b0000010111111111;
            15'd32356: log10_cal = 16'b0000010111111111;
            15'd32357: log10_cal = 16'b0000010111111111;
            15'd32358: log10_cal = 16'b0000010111111111;
            15'd32359: log10_cal = 16'b0000010111111111;
            15'd32360: log10_cal = 16'b0000010111111111;
            15'd32361: log10_cal = 16'b0000010111111111;
            15'd32362: log10_cal = 16'b0000010111111111;
            15'd32363: log10_cal = 16'b0000010111111111;
            15'd32364: log10_cal = 16'b0000010111111111;
            15'd32365: log10_cal = 16'b0000010111111111;
            15'd32366: log10_cal = 16'b0000010111111111;
            15'd32367: log10_cal = 16'b0000010111111111;
            15'd32368: log10_cal = 16'b0000010111111111;
            15'd32369: log10_cal = 16'b0000010111111111;
            15'd32370: log10_cal = 16'b0000010111111111;
            15'd32371: log10_cal = 16'b0000010111111111;
            15'd32372: log10_cal = 16'b0000010111111111;
            15'd32373: log10_cal = 16'b0000010111111111;
            15'd32374: log10_cal = 16'b0000010111111111;
            15'd32375: log10_cal = 16'b0000010111111111;
            15'd32376: log10_cal = 16'b0000010111111111;
            15'd32377: log10_cal = 16'b0000010111111111;
            15'd32378: log10_cal = 16'b0000010111111111;
            15'd32379: log10_cal = 16'b0000010111111111;
            15'd32380: log10_cal = 16'b0000010111111111;
            15'd32381: log10_cal = 16'b0000010111111111;
            15'd32382: log10_cal = 16'b0000011000000000;
            15'd32383: log10_cal = 16'b0000011000000000;
            15'd32384: log10_cal = 16'b0000011000000000;
            15'd32385: log10_cal = 16'b0000011000000000;
            15'd32386: log10_cal = 16'b0000011000000000;
            15'd32387: log10_cal = 16'b0000011000000000;
            15'd32388: log10_cal = 16'b0000011000000000;
            15'd32389: log10_cal = 16'b0000011000000000;
            15'd32390: log10_cal = 16'b0000011000000000;
            15'd32391: log10_cal = 16'b0000011000000000;
            15'd32392: log10_cal = 16'b0000011000000000;
            15'd32393: log10_cal = 16'b0000011000000000;
            15'd32394: log10_cal = 16'b0000011000000000;
            15'd32395: log10_cal = 16'b0000011000000000;
            15'd32396: log10_cal = 16'b0000011000000000;
            15'd32397: log10_cal = 16'b0000011000000000;
            15'd32398: log10_cal = 16'b0000011000000000;
            15'd32399: log10_cal = 16'b0000011000000000;
            15'd32400: log10_cal = 16'b0000011000000000;
            15'd32401: log10_cal = 16'b0000011000000000;
            15'd32402: log10_cal = 16'b0000011000000000;
            15'd32403: log10_cal = 16'b0000011000000000;
            15'd32404: log10_cal = 16'b0000011000000000;
            15'd32405: log10_cal = 16'b0000011000000000;
            15'd32406: log10_cal = 16'b0000011000000000;
            15'd32407: log10_cal = 16'b0000011000000000;
            15'd32408: log10_cal = 16'b0000011000000000;
            15'd32409: log10_cal = 16'b0000011000000000;
            15'd32410: log10_cal = 16'b0000011000000000;
            15'd32411: log10_cal = 16'b0000011000000000;
            15'd32412: log10_cal = 16'b0000011000000000;
            15'd32413: log10_cal = 16'b0000011000000000;
            15'd32414: log10_cal = 16'b0000011000000000;
            15'd32415: log10_cal = 16'b0000011000000000;
            15'd32416: log10_cal = 16'b0000011000000000;
            15'd32417: log10_cal = 16'b0000011000000000;
            15'd32418: log10_cal = 16'b0000011000000000;
            15'd32419: log10_cal = 16'b0000011000000000;
            15'd32420: log10_cal = 16'b0000011000000000;
            15'd32421: log10_cal = 16'b0000011000000000;
            15'd32422: log10_cal = 16'b0000011000000000;
            15'd32423: log10_cal = 16'b0000011000000000;
            15'd32424: log10_cal = 16'b0000011000000000;
            15'd32425: log10_cal = 16'b0000011000000000;
            15'd32426: log10_cal = 16'b0000011000000000;
            15'd32427: log10_cal = 16'b0000011000000000;
            15'd32428: log10_cal = 16'b0000011000000000;
            15'd32429: log10_cal = 16'b0000011000000000;
            15'd32430: log10_cal = 16'b0000011000000000;
            15'd32431: log10_cal = 16'b0000011000000000;
            15'd32432: log10_cal = 16'b0000011000000000;
            15'd32433: log10_cal = 16'b0000011000000000;
            15'd32434: log10_cal = 16'b0000011000000000;
            15'd32435: log10_cal = 16'b0000011000000000;
            15'd32436: log10_cal = 16'b0000011000000000;
            15'd32437: log10_cal = 16'b0000011000000000;
            15'd32438: log10_cal = 16'b0000011000000000;
            15'd32439: log10_cal = 16'b0000011000000000;
            15'd32440: log10_cal = 16'b0000011000000000;
            15'd32441: log10_cal = 16'b0000011000000000;
            15'd32442: log10_cal = 16'b0000011000000000;
            15'd32443: log10_cal = 16'b0000011000000000;
            15'd32444: log10_cal = 16'b0000011000000000;
            15'd32445: log10_cal = 16'b0000011000000000;
            15'd32446: log10_cal = 16'b0000011000000000;
            15'd32447: log10_cal = 16'b0000011000000000;
            15'd32448: log10_cal = 16'b0000011000000000;
            15'd32449: log10_cal = 16'b0000011000000000;
            15'd32450: log10_cal = 16'b0000011000000000;
            15'd32451: log10_cal = 16'b0000011000000000;
            15'd32452: log10_cal = 16'b0000011000000000;
            15'd32453: log10_cal = 16'b0000011000000000;
            15'd32454: log10_cal = 16'b0000011000000000;
            15'd32455: log10_cal = 16'b0000011000000001;
            15'd32456: log10_cal = 16'b0000011000000001;
            15'd32457: log10_cal = 16'b0000011000000001;
            15'd32458: log10_cal = 16'b0000011000000001;
            15'd32459: log10_cal = 16'b0000011000000001;
            15'd32460: log10_cal = 16'b0000011000000001;
            15'd32461: log10_cal = 16'b0000011000000001;
            15'd32462: log10_cal = 16'b0000011000000001;
            15'd32463: log10_cal = 16'b0000011000000001;
            15'd32464: log10_cal = 16'b0000011000000001;
            15'd32465: log10_cal = 16'b0000011000000001;
            15'd32466: log10_cal = 16'b0000011000000001;
            15'd32467: log10_cal = 16'b0000011000000001;
            15'd32468: log10_cal = 16'b0000011000000001;
            15'd32469: log10_cal = 16'b0000011000000001;
            15'd32470: log10_cal = 16'b0000011000000001;
            15'd32471: log10_cal = 16'b0000011000000001;
            15'd32472: log10_cal = 16'b0000011000000001;
            15'd32473: log10_cal = 16'b0000011000000001;
            15'd32474: log10_cal = 16'b0000011000000001;
            15'd32475: log10_cal = 16'b0000011000000001;
            15'd32476: log10_cal = 16'b0000011000000001;
            15'd32477: log10_cal = 16'b0000011000000001;
            15'd32478: log10_cal = 16'b0000011000000001;
            15'd32479: log10_cal = 16'b0000011000000001;
            15'd32480: log10_cal = 16'b0000011000000001;
            15'd32481: log10_cal = 16'b0000011000000001;
            15'd32482: log10_cal = 16'b0000011000000001;
            15'd32483: log10_cal = 16'b0000011000000001;
            15'd32484: log10_cal = 16'b0000011000000001;
            15'd32485: log10_cal = 16'b0000011000000001;
            15'd32486: log10_cal = 16'b0000011000000001;
            15'd32487: log10_cal = 16'b0000011000000001;
            15'd32488: log10_cal = 16'b0000011000000001;
            15'd32489: log10_cal = 16'b0000011000000001;
            15'd32490: log10_cal = 16'b0000011000000001;
            15'd32491: log10_cal = 16'b0000011000000001;
            15'd32492: log10_cal = 16'b0000011000000001;
            15'd32493: log10_cal = 16'b0000011000000001;
            15'd32494: log10_cal = 16'b0000011000000001;
            15'd32495: log10_cal = 16'b0000011000000001;
            15'd32496: log10_cal = 16'b0000011000000001;
            15'd32497: log10_cal = 16'b0000011000000001;
            15'd32498: log10_cal = 16'b0000011000000001;
            15'd32499: log10_cal = 16'b0000011000000001;
            15'd32500: log10_cal = 16'b0000011000000001;
            15'd32501: log10_cal = 16'b0000011000000001;
            15'd32502: log10_cal = 16'b0000011000000001;
            15'd32503: log10_cal = 16'b0000011000000001;
            15'd32504: log10_cal = 16'b0000011000000001;
            15'd32505: log10_cal = 16'b0000011000000001;
            15'd32506: log10_cal = 16'b0000011000000001;
            15'd32507: log10_cal = 16'b0000011000000001;
            15'd32508: log10_cal = 16'b0000011000000001;
            15'd32509: log10_cal = 16'b0000011000000001;
            15'd32510: log10_cal = 16'b0000011000000001;
            15'd32511: log10_cal = 16'b0000011000000001;
            15'd32512: log10_cal = 16'b0000011000000001;
            15'd32513: log10_cal = 16'b0000011000000001;
            15'd32514: log10_cal = 16'b0000011000000001;
            15'd32515: log10_cal = 16'b0000011000000001;
            15'd32516: log10_cal = 16'b0000011000000001;
            15'd32517: log10_cal = 16'b0000011000000001;
            15'd32518: log10_cal = 16'b0000011000000001;
            15'd32519: log10_cal = 16'b0000011000000001;
            15'd32520: log10_cal = 16'b0000011000000001;
            15'd32521: log10_cal = 16'b0000011000000001;
            15'd32522: log10_cal = 16'b0000011000000001;
            15'd32523: log10_cal = 16'b0000011000000001;
            15'd32524: log10_cal = 16'b0000011000000001;
            15'd32525: log10_cal = 16'b0000011000000001;
            15'd32526: log10_cal = 16'b0000011000000001;
            15'd32527: log10_cal = 16'b0000011000000001;
            15'd32528: log10_cal = 16'b0000011000000010;
            15'd32529: log10_cal = 16'b0000011000000010;
            15'd32530: log10_cal = 16'b0000011000000010;
            15'd32531: log10_cal = 16'b0000011000000010;
            15'd32532: log10_cal = 16'b0000011000000010;
            15'd32533: log10_cal = 16'b0000011000000010;
            15'd32534: log10_cal = 16'b0000011000000010;
            15'd32535: log10_cal = 16'b0000011000000010;
            15'd32536: log10_cal = 16'b0000011000000010;
            15'd32537: log10_cal = 16'b0000011000000010;
            15'd32538: log10_cal = 16'b0000011000000010;
            15'd32539: log10_cal = 16'b0000011000000010;
            15'd32540: log10_cal = 16'b0000011000000010;
            15'd32541: log10_cal = 16'b0000011000000010;
            15'd32542: log10_cal = 16'b0000011000000010;
            15'd32543: log10_cal = 16'b0000011000000010;
            15'd32544: log10_cal = 16'b0000011000000010;
            15'd32545: log10_cal = 16'b0000011000000010;
            15'd32546: log10_cal = 16'b0000011000000010;
            15'd32547: log10_cal = 16'b0000011000000010;
            15'd32548: log10_cal = 16'b0000011000000010;
            15'd32549: log10_cal = 16'b0000011000000010;
            15'd32550: log10_cal = 16'b0000011000000010;
            15'd32551: log10_cal = 16'b0000011000000010;
            15'd32552: log10_cal = 16'b0000011000000010;
            15'd32553: log10_cal = 16'b0000011000000010;
            15'd32554: log10_cal = 16'b0000011000000010;
            15'd32555: log10_cal = 16'b0000011000000010;
            15'd32556: log10_cal = 16'b0000011000000010;
            15'd32557: log10_cal = 16'b0000011000000010;
            15'd32558: log10_cal = 16'b0000011000000010;
            15'd32559: log10_cal = 16'b0000011000000010;
            15'd32560: log10_cal = 16'b0000011000000010;
            15'd32561: log10_cal = 16'b0000011000000010;
            15'd32562: log10_cal = 16'b0000011000000010;
            15'd32563: log10_cal = 16'b0000011000000010;
            15'd32564: log10_cal = 16'b0000011000000010;
            15'd32565: log10_cal = 16'b0000011000000010;
            15'd32566: log10_cal = 16'b0000011000000010;
            15'd32567: log10_cal = 16'b0000011000000010;
            15'd32568: log10_cal = 16'b0000011000000010;
            15'd32569: log10_cal = 16'b0000011000000010;
            15'd32570: log10_cal = 16'b0000011000000010;
            15'd32571: log10_cal = 16'b0000011000000010;
            15'd32572: log10_cal = 16'b0000011000000010;
            15'd32573: log10_cal = 16'b0000011000000010;
            15'd32574: log10_cal = 16'b0000011000000010;
            15'd32575: log10_cal = 16'b0000011000000010;
            15'd32576: log10_cal = 16'b0000011000000010;
            15'd32577: log10_cal = 16'b0000011000000010;
            15'd32578: log10_cal = 16'b0000011000000010;
            15'd32579: log10_cal = 16'b0000011000000010;
            15'd32580: log10_cal = 16'b0000011000000010;
            15'd32581: log10_cal = 16'b0000011000000010;
            15'd32582: log10_cal = 16'b0000011000000010;
            15'd32583: log10_cal = 16'b0000011000000010;
            15'd32584: log10_cal = 16'b0000011000000010;
            15'd32585: log10_cal = 16'b0000011000000010;
            15'd32586: log10_cal = 16'b0000011000000010;
            15'd32587: log10_cal = 16'b0000011000000010;
            15'd32588: log10_cal = 16'b0000011000000010;
            15'd32589: log10_cal = 16'b0000011000000010;
            15'd32590: log10_cal = 16'b0000011000000010;
            15'd32591: log10_cal = 16'b0000011000000010;
            15'd32592: log10_cal = 16'b0000011000000010;
            15'd32593: log10_cal = 16'b0000011000000010;
            15'd32594: log10_cal = 16'b0000011000000010;
            15'd32595: log10_cal = 16'b0000011000000010;
            15'd32596: log10_cal = 16'b0000011000000010;
            15'd32597: log10_cal = 16'b0000011000000010;
            15'd32598: log10_cal = 16'b0000011000000010;
            15'd32599: log10_cal = 16'b0000011000000010;
            15'd32600: log10_cal = 16'b0000011000000010;
            15'd32601: log10_cal = 16'b0000011000000011;
            15'd32602: log10_cal = 16'b0000011000000011;
            15'd32603: log10_cal = 16'b0000011000000011;
            15'd32604: log10_cal = 16'b0000011000000011;
            15'd32605: log10_cal = 16'b0000011000000011;
            15'd32606: log10_cal = 16'b0000011000000011;
            15'd32607: log10_cal = 16'b0000011000000011;
            15'd32608: log10_cal = 16'b0000011000000011;
            15'd32609: log10_cal = 16'b0000011000000011;
            15'd32610: log10_cal = 16'b0000011000000011;
            15'd32611: log10_cal = 16'b0000011000000011;
            15'd32612: log10_cal = 16'b0000011000000011;
            15'd32613: log10_cal = 16'b0000011000000011;
            15'd32614: log10_cal = 16'b0000011000000011;
            15'd32615: log10_cal = 16'b0000011000000011;
            15'd32616: log10_cal = 16'b0000011000000011;
            15'd32617: log10_cal = 16'b0000011000000011;
            15'd32618: log10_cal = 16'b0000011000000011;
            15'd32619: log10_cal = 16'b0000011000000011;
            15'd32620: log10_cal = 16'b0000011000000011;
            15'd32621: log10_cal = 16'b0000011000000011;
            15'd32622: log10_cal = 16'b0000011000000011;
            15'd32623: log10_cal = 16'b0000011000000011;
            15'd32624: log10_cal = 16'b0000011000000011;
            15'd32625: log10_cal = 16'b0000011000000011;
            15'd32626: log10_cal = 16'b0000011000000011;
            15'd32627: log10_cal = 16'b0000011000000011;
            15'd32628: log10_cal = 16'b0000011000000011;
            15'd32629: log10_cal = 16'b0000011000000011;
            15'd32630: log10_cal = 16'b0000011000000011;
            15'd32631: log10_cal = 16'b0000011000000011;
            15'd32632: log10_cal = 16'b0000011000000011;
            15'd32633: log10_cal = 16'b0000011000000011;
            15'd32634: log10_cal = 16'b0000011000000011;
            15'd32635: log10_cal = 16'b0000011000000011;
            15'd32636: log10_cal = 16'b0000011000000011;
            15'd32637: log10_cal = 16'b0000011000000011;
            15'd32638: log10_cal = 16'b0000011000000011;
            15'd32639: log10_cal = 16'b0000011000000011;
            15'd32640: log10_cal = 16'b0000011000000011;
            15'd32641: log10_cal = 16'b0000011000000011;
            15'd32642: log10_cal = 16'b0000011000000011;
            15'd32643: log10_cal = 16'b0000011000000011;
            15'd32644: log10_cal = 16'b0000011000000011;
            15'd32645: log10_cal = 16'b0000011000000011;
            15'd32646: log10_cal = 16'b0000011000000011;
            15'd32647: log10_cal = 16'b0000011000000011;
            15'd32648: log10_cal = 16'b0000011000000011;
            15'd32649: log10_cal = 16'b0000011000000011;
            15'd32650: log10_cal = 16'b0000011000000011;
            15'd32651: log10_cal = 16'b0000011000000011;
            15'd32652: log10_cal = 16'b0000011000000011;
            15'd32653: log10_cal = 16'b0000011000000011;
            15'd32654: log10_cal = 16'b0000011000000011;
            15'd32655: log10_cal = 16'b0000011000000011;
            15'd32656: log10_cal = 16'b0000011000000011;
            15'd32657: log10_cal = 16'b0000011000000011;
            15'd32658: log10_cal = 16'b0000011000000011;
            15'd32659: log10_cal = 16'b0000011000000011;
            15'd32660: log10_cal = 16'b0000011000000011;
            15'd32661: log10_cal = 16'b0000011000000011;
            15'd32662: log10_cal = 16'b0000011000000011;
            15'd32663: log10_cal = 16'b0000011000000011;
            15'd32664: log10_cal = 16'b0000011000000011;
            15'd32665: log10_cal = 16'b0000011000000011;
            15'd32666: log10_cal = 16'b0000011000000011;
            15'd32667: log10_cal = 16'b0000011000000011;
            15'd32668: log10_cal = 16'b0000011000000011;
            15'd32669: log10_cal = 16'b0000011000000011;
            15'd32670: log10_cal = 16'b0000011000000011;
            15'd32671: log10_cal = 16'b0000011000000011;
            15'd32672: log10_cal = 16'b0000011000000011;
            15'd32673: log10_cal = 16'b0000011000000011;
            15'd32674: log10_cal = 16'b0000011000000011;
            15'd32675: log10_cal = 16'b0000011000000100;
            15'd32676: log10_cal = 16'b0000011000000100;
            15'd32677: log10_cal = 16'b0000011000000100;
            15'd32678: log10_cal = 16'b0000011000000100;
            15'd32679: log10_cal = 16'b0000011000000100;
            15'd32680: log10_cal = 16'b0000011000000100;
            15'd32681: log10_cal = 16'b0000011000000100;
            15'd32682: log10_cal = 16'b0000011000000100;
            15'd32683: log10_cal = 16'b0000011000000100;
            15'd32684: log10_cal = 16'b0000011000000100;
            15'd32685: log10_cal = 16'b0000011000000100;
            15'd32686: log10_cal = 16'b0000011000000100;
            15'd32687: log10_cal = 16'b0000011000000100;
            15'd32688: log10_cal = 16'b0000011000000100;
            15'd32689: log10_cal = 16'b0000011000000100;
            15'd32690: log10_cal = 16'b0000011000000100;
            15'd32691: log10_cal = 16'b0000011000000100;
            15'd32692: log10_cal = 16'b0000011000000100;
            15'd32693: log10_cal = 16'b0000011000000100;
            15'd32694: log10_cal = 16'b0000011000000100;
            15'd32695: log10_cal = 16'b0000011000000100;
            15'd32696: log10_cal = 16'b0000011000000100;
            15'd32697: log10_cal = 16'b0000011000000100;
            15'd32698: log10_cal = 16'b0000011000000100;
            15'd32699: log10_cal = 16'b0000011000000100;
            15'd32700: log10_cal = 16'b0000011000000100;
            15'd32701: log10_cal = 16'b0000011000000100;
            15'd32702: log10_cal = 16'b0000011000000100;
            15'd32703: log10_cal = 16'b0000011000000100;
            15'd32704: log10_cal = 16'b0000011000000100;
            15'd32705: log10_cal = 16'b0000011000000100;
            15'd32706: log10_cal = 16'b0000011000000100;
            15'd32707: log10_cal = 16'b0000011000000100;
            15'd32708: log10_cal = 16'b0000011000000100;
            15'd32709: log10_cal = 16'b0000011000000100;
            15'd32710: log10_cal = 16'b0000011000000100;
            15'd32711: log10_cal = 16'b0000011000000100;
            15'd32712: log10_cal = 16'b0000011000000100;
            15'd32713: log10_cal = 16'b0000011000000100;
            15'd32714: log10_cal = 16'b0000011000000100;
            15'd32715: log10_cal = 16'b0000011000000100;
            15'd32716: log10_cal = 16'b0000011000000100;
            15'd32717: log10_cal = 16'b0000011000000100;
            15'd32718: log10_cal = 16'b0000011000000100;
            15'd32719: log10_cal = 16'b0000011000000100;
            15'd32720: log10_cal = 16'b0000011000000100;
            15'd32721: log10_cal = 16'b0000011000000100;
            15'd32722: log10_cal = 16'b0000011000000100;
            15'd32723: log10_cal = 16'b0000011000000100;
            15'd32724: log10_cal = 16'b0000011000000100;
            15'd32725: log10_cal = 16'b0000011000000100;
            15'd32726: log10_cal = 16'b0000011000000100;
            15'd32727: log10_cal = 16'b0000011000000100;
            15'd32728: log10_cal = 16'b0000011000000100;
            15'd32729: log10_cal = 16'b0000011000000100;
            15'd32730: log10_cal = 16'b0000011000000100;
            15'd32731: log10_cal = 16'b0000011000000100;
            15'd32732: log10_cal = 16'b0000011000000100;
            15'd32733: log10_cal = 16'b0000011000000100;
            15'd32734: log10_cal = 16'b0000011000000100;
            15'd32735: log10_cal = 16'b0000011000000100;
            15'd32736: log10_cal = 16'b0000011000000100;
            15'd32737: log10_cal = 16'b0000011000000100;
            15'd32738: log10_cal = 16'b0000011000000100;
            15'd32739: log10_cal = 16'b0000011000000100;
            15'd32740: log10_cal = 16'b0000011000000100;
            15'd32741: log10_cal = 16'b0000011000000100;
            15'd32742: log10_cal = 16'b0000011000000100;
            15'd32743: log10_cal = 16'b0000011000000100;
            15'd32744: log10_cal = 16'b0000011000000100;
            15'd32745: log10_cal = 16'b0000011000000100;
            15'd32746: log10_cal = 16'b0000011000000100;
            15'd32747: log10_cal = 16'b0000011000000100;
            15'd32748: log10_cal = 16'b0000011000000101;
            15'd32749: log10_cal = 16'b0000011000000101;
            15'd32750: log10_cal = 16'b0000011000000101;
            15'd32751: log10_cal = 16'b0000011000000101;
            15'd32752: log10_cal = 16'b0000011000000101;
            15'd32753: log10_cal = 16'b0000011000000101;
            15'd32754: log10_cal = 16'b0000011000000101;
            15'd32755: log10_cal = 16'b0000011000000101;
            15'd32756: log10_cal = 16'b0000011000000101;
            15'd32757: log10_cal = 16'b0000011000000101;
            15'd32758: log10_cal = 16'b0000011000000101;
            15'd32759: log10_cal = 16'b0000011000000101;
            15'd32760: log10_cal = 16'b0000011000000101;
            15'd32761: log10_cal = 16'b0000011000000101;
            15'd32762: log10_cal = 16'b0000011000000101;
            15'd32763: log10_cal = 16'b0000011000000101;
            15'd32764: log10_cal = 16'b0000011000000101;
            15'd32765: log10_cal = 16'b0000011000000101;
            15'd32766: log10_cal = 16'b0000011000000101;
            15'd32767: log10_cal = 16'b0000011000000101;
            default: log10_cal = 16'd0;
        endcase
        logtablefinish = 1'b1;
    end
    else begin
        log10_cal = 16'd0;
        logtablefinish = 1'b0;
    end
end

//log10_result
always@(posedge clk or negedge reset) begin
    if(!reset)
        log10_result <= 16'd0;
    else begin
        if(melfinish == 1'b1)
            log10_result <= log10_cal;
        else
            log10_result <= log10_result;
    end
end

//mfscoutCount
always@(posedge clk or negedge reset) begin
    if(!reset) begin
        mfscoutCount <= 6'd0;
    end
    else begin
        case(CS)
            Melcal: mfscoutCount <= mfscoutCount;
            Logtable: begin
                if(melfinish == 1'b1)
                    mfscoutCount <= mfscoutCount + 6'd1;
                else
                    mfscoutCount <= mfscoutCount;   
            end
            mfscout: mfscoutCount <= mfscoutCount;
            waitram: mfscoutCount <= mfscoutCount;
            default: mfscoutCount <= 6'd0;
        endcase
    end
end

endmodule

//fft
module fft_modulus(
    input clk,
    input div_clk,
    input reset,
    input [15:0]mixed_signal,
    input fft_s_axis_data_tvalid,
    input fft_s_axis_data_tlast,
    output fft_s_axis_data_tready,
    output fft_m_axis_data_tvalid,
    output reg modulus_done,
    output reg [15:0]result);
reg [7:0] s_axis_config_tdata;
reg s_axis_config_tvalid;
wire s_axis_config_tready;
wire [7:0] fft_m_axis_status_tdata;
wire fft_m_axis_status_tvalid;
wire fft_m_axis_data_tlast;
reg fft_m_axis_status_tready;
// OVFLO: 1bit, BLK_EXP: 8bits, XK_INDEX = 10bits
wire [7:0] m_axis_data_tuser;

wire fft_event_frame_started;
wire fft_event_tlast_unexpected;
wire fft_event_tlast_missing;
wire fft_event_status_channel_halt;
wire fft_event_data_in_channel_halt;
wire fft_event_data_out_channel_halt;

always@(posedge clk or negedge reset) begin
    if(!reset) begin
        s_axis_config_tdata <= 8'd0;
        s_axis_config_tvalid <= 1'b1;
        fft_m_axis_status_tready <= 1'b0;
    end
    else begin
        s_axis_config_tvalid <= s_axis_config_tvalid;
        if(s_axis_config_tready)
            //FWD_INV = 1, NFFT = 01010, cyclic prefix = 0, scale schedule = 0101_01010101_01010110 
            //s_axis_config_tdata <= 48'b00000101_01010101_01010110_00000001_00000000_00001010;
            s_axis_config_tdata <= 8'd0;
        else
            s_axis_config_tdata <= s_axis_config_tdata;
        if(fft_m_axis_status_tvalid)
            fft_m_axis_status_tready <= 1'b1;
        else
            fft_m_axis_status_tready <= 1'b0;
    end
end

wire [31:0] after_fft_data;

(* ram_style = "block" *)(* use_dsp = "yes" *)xfft_0 U0(
 .aclk(div_clk),
 .s_axis_config_tdata(s_axis_config_tdata),
 .s_axis_config_tvalid(s_axis_config_tvalid),
 .s_axis_config_tready(s_axis_config_tready),
 
 .s_axis_data_tdata({16'd0, mixed_signal}),
 .s_axis_data_tvalid(fft_s_axis_data_tvalid),
 .s_axis_data_tready(fft_s_axis_data_tready),
 .s_axis_data_tlast(fft_s_axis_data_tlast),
 
 .m_axis_data_tdata(after_fft_data),
 .m_axis_data_tuser(m_axis_data_tuser),
 .m_axis_data_tvalid(fft_m_axis_data_tvalid),
 .m_axis_data_tready(1'b1),
 .m_axis_data_tlast(fft_m_axis_data_tlast),
 
 .m_axis_status_tdata(fft_m_axis_status_tdata),
 .m_axis_status_tvalid(fft_m_axis_status_tvalid),
 .m_axis_status_tready(fft_m_axis_status_tready),
 
 .event_frame_started(fft_event_frame_started),
 .event_tlast_unexpected(fft_event_tlast_unexpected),
 .event_tlast_missing(fft_event_tlast_missing),
 .event_status_channel_halt(fft_event_status_channel_halt),
 .event_data_in_channel_halt(fft_event_data_in_channel_halt),
 .event_data_out_channel_halt(fft_event_data_out_channel_halt)
 );
 

wire [32:0]sum = (after_fft_data[15] == 1'b1 && after_fft_data[31] == 1'b1) ? { 17'd131071, after_fft_data[15:0]}*{ 17'd131071, after_fft_data[15:0]} + { 17'd131071, after_fft_data[31:16]}*{ 17'd131071, after_fft_data[31:16]}:
(after_fft_data[15] == 1'b1 && after_fft_data[31] == 1'b0) ? { 17'd131071, after_fft_data[15:0]}*{ 17'd131071, after_fft_data[15:0]} + { 17'd0, after_fft_data[31:16]}*{ 17'd0, after_fft_data[31:16]}:
(after_fft_data[15] == 1'b0 && after_fft_data[31] == 1'b1) ? { 17'd0, after_fft_data[15:0]}*{ 17'd0, after_fft_data[15:0]} + { 17'd131071, after_fft_data[31:16]}*{ 17'd131071, after_fft_data[31:16]}:
                                         { 17'd0, after_fft_data[15:0]}*{ 17'd0, after_fft_data[15:0]} + { 17'd0, after_fft_data[31:16]}*{ 17'd0, after_fft_data[31:16]};
 
 always@(posedge div_clk or negedge reset) begin
    if(!reset) begin
        result <= 16'b0000_0000_0000_0000;
        modulus_done <= 1'b0;
    end
    else begin
        if(!fft_m_axis_data_tvalid) begin
            result <= 16'b0000_0000_0000_0000;
            modulus_done <= 1'b0;
        end
        else begin
            result <= {sum[32], 4'b0000, sum[31:21]};
            modulus_done <= 1'b1;
        end
    end
 end
endmodule
